magic
tech sky130A
magscale 1 2
timestamp 1714754970
<< metal1 >>
rect 2848 1767 2920 2206
rect 4076 2064 4262 44152
rect 4076 1878 4104 2064
rect 4262 1878 4268 2064
rect 5418 1767 5492 2198
rect 2529 1693 2535 1767
rect 2609 1693 5492 1767
<< via1 >>
rect 4104 1878 4262 2064
rect 2535 1693 2609 1767
<< metal2 >>
rect 3416 1978 3564 2278
rect 4104 2064 4262 2070
rect 2535 1767 2609 1773
rect 2526 1693 2535 1767
rect 2609 1693 2618 1767
rect 2535 1687 2609 1693
rect 3420 964 3561 1978
rect 4095 1878 4104 2064
rect 4262 1878 4271 2064
rect 4104 1872 4262 1878
rect 4774 1244 4922 2280
rect 4774 1100 30696 1244
rect 30840 1100 30849 1244
rect 4774 1098 4922 1100
rect 3420 825 23926 964
rect 24065 825 24074 964
rect 3420 824 3561 825
<< via2 >>
rect 2535 1693 2609 1767
rect 4104 1878 4262 2064
rect 30696 1100 30840 1244
rect 23926 825 24065 964
<< metal3 >>
rect 4099 2064 4109 2069
rect 4099 1878 4104 2064
rect 4099 1873 4109 1878
rect 4267 1873 4273 2069
rect 2516 1772 2632 1788
rect 2516 1688 2530 1772
rect 2604 1767 2632 1772
rect 2609 1693 2632 1767
rect 2604 1688 2632 1693
rect 2516 1658 2632 1688
rect 30691 1244 30701 1249
rect 30691 1100 30696 1244
rect 30691 1095 30701 1100
rect 30845 1095 30851 1249
rect 23921 964 23931 969
rect 23921 825 23926 964
rect 23921 820 23931 825
rect 24070 820 24076 969
<< via3 >>
rect 4109 2064 4267 2069
rect 4109 1878 4262 2064
rect 4262 1878 4267 2064
rect 4109 1873 4267 1878
rect 2530 1767 2604 1772
rect 2530 1693 2535 1767
rect 2535 1693 2604 1767
rect 2530 1688 2604 1693
rect 30701 1244 30845 1249
rect 30701 1100 30840 1244
rect 30840 1100 30845 1244
rect 30701 1095 30845 1100
rect 23931 964 24070 969
rect 23931 825 24065 964
rect 24065 825 24070 964
rect 23931 820 24070 825
<< metal4 >>
rect 798 44616 858 45152
rect 1534 44616 1594 45152
rect 2270 44616 2330 45152
rect 3006 44616 3066 45152
rect 3742 44616 3802 45152
rect 4478 44616 4538 45152
rect 5214 44616 5274 45152
rect 5950 44616 6010 45152
rect 6686 44616 6746 45152
rect 7422 44616 7482 45152
rect 8158 44616 8218 45152
rect 8894 44616 8954 45152
rect 9630 44616 9690 45152
rect 10366 44616 10426 45152
rect 11102 44616 11162 45152
rect 11838 44616 11898 45152
rect 12574 44616 12634 45152
rect 13310 44616 13370 45152
rect 14046 44616 14106 45152
rect 14782 44616 14842 45152
rect 15518 44616 15578 45152
rect 16254 44616 16314 45152
rect 16990 44616 17050 45152
rect 17726 44616 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 172 44298 31790 44616
rect 200 1778 500 44152
rect 4108 2069 4268 2070
rect 4108 1873 4109 2069
rect 4267 2050 4268 2069
rect 9800 2050 10100 44298
rect 4267 1892 10100 2050
rect 4267 1873 4268 1892
rect 4108 1872 4268 1873
rect 200 1770 1378 1778
rect 2529 1772 2605 1773
rect 200 1767 1592 1770
rect 2529 1767 2530 1772
rect 200 1693 2530 1767
rect 200 1691 1592 1693
rect 200 1683 1378 1691
rect 2529 1688 2530 1693
rect 2604 1688 2605 1772
rect 2529 1687 2605 1688
rect 200 1000 500 1683
rect 9800 1000 10100 1892
rect 30700 1249 30846 1250
rect 30700 1095 30701 1249
rect 30845 1244 30846 1249
rect 30845 1100 31408 1244
rect 30845 1095 30846 1100
rect 30700 1094 30846 1095
rect 23930 969 24071 970
rect 23930 820 23931 969
rect 24070 964 24071 969
rect 24070 825 27021 964
rect 24070 820 24071 825
rect 23930 819 24071 820
rect 26882 200 27021 825
rect 31264 200 31408 1100
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31264 112 31462 200
rect 31282 0 31462 112
use oscillator_20MHZ  oscillator_20MHZ_0
timestamp 1714689377
transform 0 1 3590 -1 0 43760
box -396 600 41608 1900
use oscillator_21MHZ  oscillator_21MHZ_0
timestamp 1714689377
transform 0 -1 4750 -1 0 44148
box 4 600 41996 1900
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
