magic
tech sky130A
magscale 1 2
timestamp 1716504190
<< pwell >>
rect -361 -2596 361 2596
<< psubdiff >>
rect -325 2526 -229 2560
rect 229 2526 325 2560
rect -325 2464 -291 2526
rect 291 2464 325 2526
rect -325 -2526 -291 -2464
rect 291 -2526 325 -2464
rect -325 -2560 -229 -2526
rect 229 -2560 325 -2526
<< psubdiffcont >>
rect -229 2526 229 2560
rect -325 -2464 -291 2464
rect 291 -2464 325 2464
rect -229 -2560 229 -2526
<< poly >>
rect -195 2414 -129 2430
rect -195 2380 -179 2414
rect -145 2380 -129 2414
rect -195 2000 -129 2380
rect -195 -2380 -129 -2000
rect -195 -2414 -179 -2380
rect -145 -2414 -129 -2380
rect -195 -2430 -129 -2414
rect -87 2414 -21 2430
rect -87 2380 -71 2414
rect -37 2380 -21 2414
rect -87 2000 -21 2380
rect -87 -2380 -21 -2000
rect -87 -2414 -71 -2380
rect -37 -2414 -21 -2380
rect -87 -2430 -21 -2414
rect 21 2414 87 2430
rect 21 2380 37 2414
rect 71 2380 87 2414
rect 21 2000 87 2380
rect 21 -2380 87 -2000
rect 21 -2414 37 -2380
rect 71 -2414 87 -2380
rect 21 -2430 87 -2414
rect 129 2414 195 2430
rect 129 2380 145 2414
rect 179 2380 195 2414
rect 129 2000 195 2380
rect 129 -2380 195 -2000
rect 129 -2414 145 -2380
rect 179 -2414 195 -2380
rect 129 -2430 195 -2414
<< polycont >>
rect -179 2380 -145 2414
rect -179 -2414 -145 -2380
rect -71 2380 -37 2414
rect -71 -2414 -37 -2380
rect 37 2380 71 2414
rect 37 -2414 71 -2380
rect 145 2380 179 2414
rect 145 -2414 179 -2380
<< npolyres >>
rect -195 -2000 -129 2000
rect -87 -2000 -21 2000
rect 21 -2000 87 2000
rect 129 -2000 195 2000
<< locali >>
rect -325 2526 -229 2560
rect 229 2526 325 2560
rect -325 2464 -291 2526
rect 291 2464 325 2526
rect -195 2380 -179 2414
rect -145 2380 -129 2414
rect -87 2380 -71 2414
rect -37 2380 -21 2414
rect 21 2380 37 2414
rect 71 2380 87 2414
rect 129 2380 145 2414
rect 179 2380 195 2414
rect -195 -2414 -179 -2380
rect -145 -2414 -129 -2380
rect -87 -2414 -71 -2380
rect -37 -2414 -21 -2380
rect 21 -2414 37 -2380
rect 71 -2414 87 -2380
rect 129 -2414 145 -2380
rect 179 -2414 195 -2380
rect -325 -2526 -291 -2464
rect 291 -2526 325 -2464
rect -325 -2560 -229 -2526
rect 229 -2560 325 -2526
<< viali >>
rect -179 2380 -145 2414
rect -71 2380 -37 2414
rect 37 2380 71 2414
rect 145 2380 179 2414
rect -179 2017 -145 2380
rect -71 2017 -37 2380
rect 37 2017 71 2380
rect 145 2017 179 2380
rect -179 -2380 -145 -2017
rect -71 -2380 -37 -2017
rect 37 -2380 71 -2017
rect 145 -2380 179 -2017
rect -179 -2414 -145 -2380
rect -71 -2414 -37 -2380
rect 37 -2414 71 -2380
rect 145 -2414 179 -2380
<< metal1 >>
rect -185 2414 -139 2426
rect -185 2017 -179 2414
rect -145 2017 -139 2414
rect -185 2005 -139 2017
rect -77 2414 -31 2426
rect -77 2017 -71 2414
rect -37 2017 -31 2414
rect -77 2005 -31 2017
rect 31 2414 77 2426
rect 31 2017 37 2414
rect 71 2017 77 2414
rect 31 2005 77 2017
rect 139 2414 185 2426
rect 139 2017 145 2414
rect 179 2017 185 2414
rect 139 2005 185 2017
rect -185 -2017 -139 -2005
rect -185 -2414 -179 -2017
rect -145 -2414 -139 -2017
rect -185 -2426 -139 -2414
rect -77 -2017 -31 -2005
rect -77 -2414 -71 -2017
rect -37 -2414 -31 -2017
rect -77 -2426 -31 -2414
rect 31 -2017 77 -2005
rect 31 -2414 37 -2017
rect 71 -2414 77 -2017
rect 31 -2426 77 -2414
rect 139 -2017 185 -2005
rect 139 -2414 145 -2017
rect 179 -2414 185 -2017
rect 139 -2426 185 -2414
<< properties >>
string FIXED_BBOX -308 -2543 308 2543
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.330 l 20 m 1 nx 4 wmin 0.330 lmin 1.650 rho 48.2 val 2.921k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
