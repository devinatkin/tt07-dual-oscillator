magic
tech sky130A
timestamp 1715222833
<< nwell >>
rect 451 1212 914 1657
<< pwell >>
rect 451 834 914 1212
<< psubdiff >>
rect 469 1178 512 1195
rect 558 1178 608 1195
rect 763 1178 805 1195
rect 851 1178 892 1195
rect 469 1162 486 1178
rect 469 862 486 885
rect 875 862 892 1178
rect 469 845 510 862
rect 567 845 596 862
rect 777 845 805 862
rect 857 845 892 862
<< nsubdiff >>
rect 469 1622 499 1639
rect 848 1622 896 1639
rect 469 1609 486 1622
rect 469 1247 486 1266
rect 875 1247 896 1622
rect 469 1230 499 1247
rect 866 1230 896 1247
<< psubdiffcont >>
rect 512 1178 558 1195
rect 805 1178 851 1195
rect 469 885 486 1162
rect 510 845 567 862
rect 805 845 857 862
<< nsubdiffcont >>
rect 499 1622 848 1639
rect 469 1266 486 1609
rect 499 1230 866 1247
<< locali >>
rect 469 1622 499 1640
rect 866 1622 896 1640
rect 469 1609 486 1622
rect 468 1266 469 1321
rect 468 1247 486 1266
rect 875 1247 896 1622
rect 468 1241 499 1247
rect 469 1230 499 1241
rect 866 1230 896 1247
rect 469 1178 512 1195
rect 558 1178 805 1195
rect 851 1178 896 1195
rect 469 1162 487 1178
rect 486 885 487 1162
rect 469 862 487 885
rect 875 862 896 1178
rect 469 845 486 862
rect 597 845 805 862
rect 862 845 896 862
<< viali >>
rect 499 1639 866 1640
rect 499 1622 848 1639
rect 848 1622 866 1639
rect 486 845 510 862
rect 510 845 567 862
rect 567 845 597 862
rect 818 845 857 862
rect 857 845 862 862
rect 486 844 597 845
<< metal1 >>
rect 451 1640 914 1657
rect 451 1622 499 1640
rect 866 1622 914 1640
rect 451 1609 914 1622
rect 451 1586 875 1609
rect 451 1567 689 1586
rect 734 1567 875 1586
rect 893 1567 914 1609
rect 566 1479 605 1531
rect 655 1479 832 1531
rect 551 1398 568 1413
rect 551 1346 832 1398
rect 551 1247 568 1346
rect 473 1178 568 1247
rect 551 1123 568 1178
rect 590 1247 794 1316
rect 835 1247 897 1248
rect 590 1178 897 1247
rect 590 1144 794 1178
rect 551 1105 616 1123
rect 551 1053 772 1105
rect 551 1039 616 1053
rect 598 926 687 978
rect 735 926 771 978
rect 800 889 914 890
rect 788 888 914 889
rect 451 884 914 888
rect 451 862 605 884
rect 451 844 486 862
rect 597 844 605 862
rect 451 839 605 844
rect 652 862 914 884
rect 652 845 818 862
rect 862 845 914 862
rect 652 839 914 845
rect 451 834 914 839
<< via1 >>
rect 689 1559 734 1586
rect 605 1479 655 1531
rect 687 926 735 978
rect 605 839 652 884
<< metal2 >>
rect 682 1586 739 1590
rect 682 1559 689 1586
rect 734 1559 739 1586
rect 601 1531 658 1535
rect 601 1479 605 1531
rect 655 1479 658 1531
rect 601 884 658 1479
rect 682 978 739 1559
rect 682 926 687 978
rect 735 926 739 978
rect 682 920 739 926
rect 601 839 605 884
rect 652 839 658 884
rect 601 836 658 839
use sky130_fd_pr__nfet_01v8_EEHCG5  sky130_fd_pr__nfet_01v8_EEHCG5_0
timestamp 1715222833
transform 0 -1 685 1 0 1081
box -79 -94 79 94
use sky130_fd_pr__nfet_01v8_EEHCG5  sky130_fd_pr__nfet_01v8_EEHCG5_1
timestamp 1715222833
transform 0 -1 685 1 0 952
box -79 -94 79 94
use sky130_fd_pr__pfet_01v8_BPT9FA  sky130_fd_pr__pfet_01v8_BPT9FA_0
timestamp 1715222833
transform 0 -1 692 1 0 1371
box -97 -150 97 150
use sky130_fd_pr__pfet_01v8_BPT9FA  XM3
timestamp 1715222833
transform 0 -1 692 1 0 1500
box -97 -150 97 150
<< labels >>
flabel metal1 473 1178 558 1247 0 FreeSans 400 0 0 0 IN
port 0 nsew
flabel metal1 590 1178 879 1247 0 FreeSans 400 0 0 0 OUT
port 1 nsew
flabel metal1 451 1567 499 1657 0 FreeSans 400 0 0 0 VCC
port 2 nsew
flabel metal1 451 834 486 888 0 FreeSans 400 0 0 0 VSS
port 4 nsew
<< end >>
