magic
tech sky130A
timestamp 1716849570
<< nwell >>
rect 0 0 1387 1710
<< nsubdiff >>
rect 42 1627 92 1645
rect 1279 1627 1344 1645
rect 42 1598 60 1627
rect 42 52 60 68
rect 1326 1592 1344 1627
rect 1326 52 1344 62
rect 42 34 100 52
rect 1287 34 1344 52
<< nsubdiffcont >>
rect 92 1627 1279 1645
rect 42 68 60 1598
rect 1326 62 1344 1592
rect 100 34 1287 52
<< locali >>
rect 42 1627 92 1645
rect 1279 1627 1344 1645
rect 42 1598 60 1627
rect 42 52 60 68
rect 1326 1592 1344 1627
rect 1326 52 1344 62
rect 42 34 100 52
rect 1287 34 1344 52
<< viali >>
rect 103 1627 1270 1645
rect 42 727 60 789
rect 1326 716 1344 822
<< metal1 >>
rect 42 1669 1344 1677
rect 42 1629 101 1669
rect 178 1645 1344 1669
rect 42 1627 103 1629
rect 1270 1627 1344 1645
rect 42 1621 1344 1627
rect 141 1599 1093 1602
rect 141 1572 263 1599
rect 311 1572 1121 1599
rect 141 1569 1121 1572
rect 202 1518 228 1569
rect 1084 1527 1121 1569
rect 113 1143 157 1148
rect 113 1053 120 1143
rect 150 1053 157 1143
rect 552 1139 599 1146
rect 195 1032 224 1128
rect 552 1060 557 1139
rect 592 1060 599 1139
rect 552 1052 599 1060
rect 640 1129 712 1146
rect 640 1055 653 1129
rect 699 1055 712 1129
rect 640 1049 712 1055
rect 1006 1136 1052 1146
rect 1006 1057 1011 1136
rect 1042 1057 1052 1136
rect 1006 1046 1052 1057
rect 1090 1032 1125 1129
rect 146 1030 1125 1032
rect 146 1003 266 1030
rect 314 1004 1125 1030
rect 314 1003 1098 1004
rect 146 999 1098 1003
rect 88 975 1134 980
rect 88 946 118 975
rect 146 974 1134 975
rect 146 946 563 974
rect 88 945 563 946
rect 591 945 1134 974
rect 88 941 1134 945
rect 93 880 1142 887
rect 93 833 188 880
rect 225 879 1142 880
rect 225 833 638 879
rect 694 878 1142 879
rect 694 833 1087 878
rect 93 829 1087 833
rect 1133 829 1142 878
rect 93 823 1142 829
rect 1308 822 1357 831
rect 27 789 75 792
rect 27 727 42 789
rect 60 775 75 789
rect 1308 775 1326 822
rect 60 770 1326 775
rect 60 769 1021 770
rect 60 740 119 769
rect 147 740 572 769
rect 600 741 1021 769
rect 1049 741 1326 770
rect 600 740 1326 741
rect 60 736 1326 740
rect 60 727 75 736
rect 27 724 75 727
rect 1308 716 1326 736
rect 1344 716 1357 822
rect 1308 708 1357 716
rect 143 700 1095 704
rect 143 673 266 700
rect 314 673 1095 700
rect 143 671 1095 673
rect 194 648 244 654
rect 101 630 158 636
rect 101 573 114 630
rect 150 573 158 630
rect 194 598 202 648
rect 238 598 244 648
rect 194 592 244 598
rect 559 632 616 641
rect 101 564 158 573
rect 559 575 564 632
rect 610 575 616 632
rect 559 569 616 575
rect 661 572 696 671
rect 1098 650 1145 653
rect 1004 641 1054 647
rect 1004 572 1008 641
rect 1047 572 1054 641
rect 1098 592 1104 650
rect 1140 592 1145 650
rect 1098 587 1145 592
rect 1004 565 1054 572
rect 653 134 678 167
rect 144 132 1096 134
rect 144 105 264 132
rect 312 105 1096 132
rect 144 101 1096 105
<< via1 >>
rect 101 1645 178 1669
rect 101 1629 103 1645
rect 103 1629 178 1645
rect 263 1572 311 1599
rect 120 1053 150 1143
rect 557 1060 592 1139
rect 653 1055 699 1129
rect 1011 1057 1042 1136
rect 266 1003 314 1030
rect 118 946 146 975
rect 563 945 591 974
rect 188 833 225 880
rect 638 833 694 879
rect 1087 829 1133 878
rect 119 740 147 769
rect 572 740 600 769
rect 1021 741 1049 770
rect 266 673 314 700
rect 114 573 150 630
rect 202 598 238 648
rect 564 575 610 632
rect 1008 572 1047 641
rect 1104 592 1140 650
rect 264 105 312 132
<< metal2 >>
rect 110 1677 162 1678
rect 93 1669 189 1677
rect 93 1629 101 1669
rect 178 1629 189 1669
rect 93 1622 189 1629
rect 110 1143 162 1622
rect 110 1053 120 1143
rect 150 1053 162 1143
rect 110 1048 162 1053
rect 257 1599 321 1602
rect 257 1572 263 1599
rect 311 1572 321 1599
rect 110 1044 155 1048
rect 113 982 150 1044
rect 257 1030 321 1572
rect 552 1139 599 1146
rect 552 1060 557 1139
rect 592 1060 599 1139
rect 640 1129 712 1146
rect 640 1121 653 1129
rect 552 1052 599 1060
rect 639 1055 653 1121
rect 699 1055 712 1129
rect 257 1003 266 1030
rect 314 1003 321 1030
rect 112 975 152 982
rect 112 946 118 975
rect 146 946 152 975
rect 112 769 152 946
rect 167 880 243 891
rect 167 833 188 880
rect 225 833 243 880
rect 167 797 243 833
rect 112 740 119 769
rect 147 740 152 769
rect 112 730 152 740
rect 113 636 150 730
rect 197 655 237 797
rect 257 700 321 1003
rect 559 974 596 1052
rect 559 945 563 974
rect 591 945 596 974
rect 559 938 596 945
rect 639 1049 712 1055
rect 1006 1136 1053 1146
rect 1006 1057 1011 1136
rect 1042 1057 1053 1136
rect 563 774 594 938
rect 639 889 679 1049
rect 1006 1046 1053 1057
rect 1016 940 1053 1046
rect 627 879 707 889
rect 627 833 638 879
rect 694 833 707 879
rect 627 823 707 833
rect 1017 774 1048 940
rect 1081 878 1142 886
rect 1081 829 1087 878
rect 1133 829 1142 878
rect 1081 821 1142 829
rect 563 769 603 774
rect 563 740 572 769
rect 600 740 603 769
rect 563 739 603 740
rect 257 673 266 700
rect 314 673 321 700
rect 194 648 241 655
rect 101 630 158 636
rect 101 573 114 630
rect 150 573 158 630
rect 194 598 202 648
rect 238 598 241 648
rect 194 592 241 598
rect 101 564 158 573
rect 257 132 321 673
rect 566 641 603 739
rect 1013 770 1050 774
rect 1013 741 1021 770
rect 1049 741 1050 770
rect 1013 647 1050 741
rect 1097 653 1137 821
rect 1097 650 1145 653
rect 1004 641 1054 647
rect 559 632 616 641
rect 559 575 564 632
rect 610 575 616 632
rect 559 569 616 575
rect 1004 572 1008 641
rect 1047 572 1054 641
rect 1097 592 1104 650
rect 1140 592 1145 650
rect 1097 589 1145 592
rect 1098 587 1145 589
rect 566 568 603 569
rect 1004 565 1054 572
rect 257 105 264 132
rect 312 105 321 132
rect 257 102 321 105
use sky130_fd_pr__pfet_01v8_lvt_NFH92T  sky130_fd_pr__pfet_01v8_lvt_NFH92T_0
timestamp 1716849570
transform 1 0 622 0 1 1300
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_0
timestamp 1716849570
transform 1 0 1072 0 1 1300
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_1
timestamp 1716849570
transform 1 0 172 0 1 1300
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_2
timestamp 1716849570
transform 1 0 172 0 1 400
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_3
timestamp 1716849570
transform 1 0 622 0 1 400
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_4
timestamp 1716849570
transform 1 0 1072 0 1 400
box -72 -300 72 300
<< labels >>
flabel metal2 225 823 232 825 0 FreeSans 240 0 0 0 DB
port 4 nsew
flabel metal1 312 101 1096 134 0 FreeSans 240 0 0 0 DA
port 5 nsew
flabel metal1 147 736 572 775 0 FreeSans 240 0 0 0 VCC
port 6 nsew
<< end >>
