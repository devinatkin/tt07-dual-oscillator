magic
tech sky130A
timestamp 1717178954
<< nwell >>
rect -114 738 1613 1473
<< pwell >>
rect -114 -82 1613 738
<< psubdiff >>
rect -68 662 -22 679
rect 1502 662 1581 679
rect -68 617 -50 662
rect -68 -35 -50 -19
rect 1563 630 1581 662
rect 1563 -35 1581 -16
rect -68 -52 -21 -35
rect 1503 -52 1581 -35
<< nsubdiff >>
rect -68 1420 -7 1437
rect 1165 1420 1242 1437
rect -68 1373 -51 1420
rect -68 777 -51 800
rect 1225 1371 1242 1420
rect 1225 777 1242 798
rect -68 760 -22 777
rect 1150 760 1242 777
<< psubdiffcont >>
rect -22 662 1502 679
rect -68 -19 -50 617
rect 1563 -16 1581 630
rect -21 -52 1503 -35
<< nsubdiffcont >>
rect -7 1420 1165 1437
rect -68 800 -51 1373
rect 1225 798 1242 1371
rect -22 760 1150 777
<< locali >>
rect -68 1420 -7 1437
rect 1165 1420 1242 1437
rect -68 1373 -51 1420
rect -68 777 -51 800
rect 1225 1371 1242 1420
rect 1225 777 1242 798
rect -68 760 -22 777
rect 1150 760 1242 777
rect -68 662 -22 679
rect 1502 662 1581 679
rect -68 617 -50 662
rect -68 -35 -50 -19
rect 1563 630 1581 662
rect 1563 -35 1581 -16
rect -68 -52 -21 -35
rect 1503 -52 1581 -35
<< viali >>
rect 76 1420 190 1437
rect 300 1420 414 1437
rect 530 1420 644 1437
rect 774 1420 888 1437
rect 1014 1420 1128 1437
rect 70 -52 217 -35
rect 353 -52 500 -35
rect 588 -52 735 -35
rect 840 -52 987 -35
rect 1098 -52 1245 -35
rect 1355 -52 1502 -35
<< metal1 >>
rect -68 1449 1296 1455
rect -68 1437 381 1449
rect 521 1437 1296 1449
rect -68 1420 76 1437
rect 190 1420 300 1437
rect 521 1420 530 1437
rect 644 1420 774 1437
rect 888 1420 1014 1437
rect 1128 1420 1296 1437
rect -68 1413 1296 1420
rect 42 1369 1137 1399
rect 98 1330 133 1337
rect 98 1233 103 1330
rect 132 1233 133 1330
rect 98 1225 133 1233
rect 255 1332 289 1338
rect 567 1336 609 1342
rect 255 1234 261 1332
rect 287 1234 289 1332
rect 255 1226 289 1234
rect 413 1331 449 1335
rect 413 1231 416 1331
rect 445 1231 449 1331
rect 413 1226 449 1231
rect 567 1231 570 1336
rect 604 1231 609 1336
rect 567 1226 609 1231
rect 722 1334 768 1341
rect 722 1231 727 1334
rect 761 1231 768 1334
rect 722 1226 768 1231
rect 882 1330 924 1336
rect 882 1234 887 1330
rect 918 1234 924 1330
rect 882 1226 924 1234
rect 1039 1328 1082 1334
rect 1039 1232 1044 1328
rect 1076 1232 1082 1328
rect 1039 1226 1082 1232
rect 15 987 50 992
rect 15 874 23 987
rect 15 866 50 874
rect 171 987 207 991
rect 171 873 175 987
rect 202 873 207 987
rect 171 865 207 873
rect 330 987 366 992
rect 330 873 334 987
rect 361 873 366 987
rect 330 866 366 873
rect 490 987 526 992
rect 490 873 495 987
rect 522 873 526 987
rect 490 866 526 873
rect 650 988 684 992
rect 650 871 652 988
rect 681 871 684 988
rect 650 866 684 871
rect 803 988 837 992
rect 803 871 807 988
rect 834 871 837 988
rect 803 866 837 871
rect 966 988 1000 992
rect 966 872 970 988
rect 997 872 1000 988
rect 966 866 1000 872
rect 1124 987 1159 992
rect 1124 871 1128 987
rect 1155 871 1159 987
rect 1124 866 1159 871
rect 43 804 1139 834
rect 43 738 138 804
rect 25 593 120 645
rect 25 562 1509 593
rect 73 530 113 536
rect -3 177 31 530
rect 73 419 79 530
rect 107 419 113 530
rect 73 415 113 419
rect 236 527 272 536
rect 236 420 242 527
rect 268 420 272 527
rect 74 414 110 415
rect 236 414 272 420
rect 393 532 428 538
rect 393 419 396 532
rect 424 419 428 532
rect 393 414 428 419
rect 554 523 590 528
rect 554 419 558 523
rect 585 419 590 523
rect 554 413 590 419
rect 710 520 744 526
rect 710 419 715 520
rect 741 419 744 520
rect 710 414 744 419
rect 869 521 904 529
rect 869 419 874 521
rect 900 419 904 521
rect 869 414 904 419
rect 1026 521 1062 533
rect 1026 419 1030 521
rect 1056 419 1062 521
rect 1026 414 1062 419
rect 1185 521 1220 529
rect 1185 419 1190 521
rect 1216 419 1220 521
rect 1185 414 1220 419
rect 1336 525 1378 533
rect 1336 419 1344 525
rect 1372 419 1378 525
rect 1336 415 1378 419
rect 1501 525 1537 533
rect 1501 418 1505 525
rect 1533 418 1537 525
rect 1341 414 1375 415
rect 1501 413 1537 418
rect -3 73 0 177
rect 28 73 31 177
rect -3 46 31 73
rect 152 183 192 191
rect 152 79 159 183
rect 187 79 192 183
rect 152 63 192 79
rect 312 184 352 191
rect 312 73 319 184
rect 347 73 352 184
rect 312 63 352 73
rect 471 182 511 192
rect 471 69 476 182
rect 504 69 511 182
rect 471 59 511 69
rect 624 184 669 190
rect 624 69 634 184
rect 660 69 669 184
rect 624 64 669 69
rect 789 186 824 191
rect 789 70 794 186
rect 820 70 824 186
rect 789 65 824 70
rect 945 185 981 191
rect 945 71 949 185
rect 976 71 981 185
rect 945 64 981 71
rect 1105 187 1141 191
rect 1105 70 1111 187
rect 1137 70 1141 187
rect 1105 63 1141 70
rect 1264 186 1303 191
rect 1264 70 1270 186
rect 1298 70 1303 186
rect 1264 64 1303 70
rect 1422 186 1458 192
rect 1422 68 1425 186
rect 1454 68 1458 186
rect 1422 64 1458 68
rect 26 -4 1510 27
rect -68 -25 1581 -21
rect -68 -35 617 -25
rect 690 -35 1581 -25
rect -68 -52 70 -35
rect 217 -52 353 -35
rect 500 -52 588 -35
rect 735 -52 840 -35
rect 987 -52 1098 -35
rect 1245 -52 1355 -35
rect 1502 -52 1581 -35
rect -68 -56 617 -52
rect 690 -56 1581 -52
rect -68 -63 1581 -56
<< via1 >>
rect 381 1437 521 1449
rect 381 1420 414 1437
rect 414 1420 521 1437
rect 103 1233 132 1330
rect 261 1234 287 1332
rect 416 1231 445 1331
rect 570 1231 604 1336
rect 727 1231 761 1334
rect 887 1234 918 1330
rect 1044 1232 1076 1328
rect 23 874 50 987
rect 175 873 202 987
rect 334 873 361 987
rect 495 873 522 987
rect 652 871 681 988
rect 807 871 834 988
rect 970 872 997 988
rect 1128 871 1155 987
rect 79 419 107 530
rect 242 420 268 527
rect 396 419 424 532
rect 558 419 585 523
rect 715 419 741 520
rect 874 419 900 521
rect 1030 419 1056 521
rect 1190 419 1216 521
rect 1344 419 1372 525
rect 1505 418 1533 525
rect 0 73 28 177
rect 159 79 187 183
rect 319 73 347 184
rect 476 69 504 182
rect 634 69 660 184
rect 794 70 820 186
rect 949 71 976 185
rect 1111 70 1137 187
rect 1270 70 1298 186
rect 1425 68 1454 186
rect 617 -35 690 -25
rect 617 -52 690 -35
rect 617 -56 690 -52
<< metal2 >>
rect 370 1449 529 1456
rect 370 1420 381 1449
rect 521 1420 529 1449
rect 370 1413 529 1420
rect 16 987 50 1339
rect 98 1330 133 1337
rect 98 1233 103 1330
rect 132 1233 133 1330
rect 98 1225 133 1233
rect 16 985 23 987
rect 16 872 21 985
rect 49 872 50 874
rect 16 855 50 872
rect 99 853 133 1225
rect 172 991 206 1334
rect 255 1332 294 1340
rect 255 1234 261 1332
rect 290 1234 294 1332
rect 255 1225 294 1234
rect 171 987 207 991
rect 171 873 175 987
rect 203 873 207 987
rect 171 865 207 873
rect 172 850 206 865
rect 255 854 289 1225
rect 331 992 365 1338
rect 407 1331 455 1413
rect 407 1231 416 1331
rect 445 1231 455 1331
rect 407 1225 455 1231
rect 330 987 366 992
rect 330 873 334 987
rect 362 873 366 987
rect 330 866 366 873
rect 331 854 365 866
rect 414 850 448 1225
rect 491 992 525 1344
rect 570 1342 604 1343
rect 567 1336 609 1342
rect 567 1231 570 1336
rect 604 1231 609 1336
rect 567 1226 609 1231
rect 490 987 526 992
rect 490 945 495 987
rect 489 873 495 945
rect 523 873 526 987
rect 489 693 526 873
rect 570 859 604 1226
rect 650 988 684 1345
rect 722 1334 768 1341
rect 722 1231 727 1334
rect 761 1231 768 1334
rect 722 1226 768 1231
rect 650 871 652 988
rect 681 871 684 988
rect 650 861 684 871
rect 726 857 760 1226
rect 803 988 837 1339
rect 882 1330 924 1336
rect 882 1234 887 1330
rect 918 1234 924 1330
rect 882 1226 924 1234
rect 803 871 807 988
rect 836 871 837 988
rect 803 855 837 871
rect 886 848 920 1226
rect 966 988 1000 1333
rect 1039 1328 1082 1334
rect 1039 1232 1044 1328
rect 1076 1232 1082 1328
rect 1039 1226 1082 1232
rect 966 872 970 988
rect 998 872 1000 988
rect 966 849 1000 872
rect 1043 849 1077 1226
rect 1125 992 1159 1335
rect 1124 987 1159 992
rect 1124 871 1128 987
rect 1156 871 1159 987
rect 1124 866 1159 871
rect 1125 851 1159 866
rect 487 660 593 693
rect 73 530 113 536
rect -3 177 31 530
rect 73 419 79 530
rect 107 419 113 530
rect 73 415 113 419
rect -3 73 0 177
rect 28 73 31 177
rect -3 46 31 73
rect 75 50 109 415
rect 154 183 188 539
rect 154 79 159 183
rect 187 79 188 183
rect 154 55 188 79
rect 237 527 271 536
rect 237 420 242 527
rect 270 420 271 527
rect 237 52 271 420
rect 314 191 348 541
rect 393 532 428 538
rect 393 419 396 532
rect 424 419 428 532
rect 393 414 428 419
rect 312 184 352 191
rect 312 73 319 184
rect 347 73 352 184
rect 312 63 352 73
rect 314 57 348 63
rect 394 54 428 414
rect 474 182 508 533
rect 554 523 591 660
rect 554 419 558 523
rect 587 420 591 523
rect 587 419 590 420
rect 554 413 590 419
rect 474 69 476 182
rect 504 69 508 182
rect 474 49 508 69
rect 555 44 589 413
rect 630 191 664 528
rect 710 520 744 526
rect 710 419 715 520
rect 623 185 669 191
rect 623 69 634 185
rect 664 69 669 185
rect 623 -21 669 69
rect 710 42 744 419
rect 789 186 823 529
rect 869 521 904 529
rect 869 419 874 521
rect 902 419 904 521
rect 869 414 904 419
rect 789 70 794 186
rect 822 70 823 186
rect 789 45 823 70
rect 870 45 904 414
rect 946 186 980 534
rect 1026 521 1062 533
rect 1026 419 1030 521
rect 1058 419 1062 521
rect 1026 414 1062 419
rect 946 71 949 186
rect 978 71 980 186
rect 946 50 980 71
rect 1027 49 1061 414
rect 1106 187 1140 531
rect 1106 70 1111 187
rect 1139 70 1140 187
rect 1106 47 1140 70
rect 1185 521 1220 529
rect 1185 419 1190 521
rect 1218 419 1220 521
rect 1185 414 1220 419
rect 1185 45 1219 414
rect 1265 191 1299 528
rect 1336 525 1378 533
rect 1336 419 1344 525
rect 1372 419 1378 525
rect 1336 415 1378 419
rect 1264 186 1303 191
rect 1264 70 1270 186
rect 1298 70 1303 186
rect 1264 64 1303 70
rect 1265 44 1299 64
rect 1341 45 1375 415
rect 1423 192 1457 529
rect 1501 525 1537 533
rect 1501 418 1505 525
rect 1533 418 1537 525
rect 1501 413 1537 418
rect 1422 186 1458 192
rect 1422 68 1425 186
rect 1454 68 1458 186
rect 1422 64 1458 68
rect 1423 45 1457 64
rect 1502 44 1536 413
rect 609 -25 695 -21
rect 609 -56 617 -25
rect 690 -56 695 -25
rect 609 -63 695 -56
<< via2 >>
rect 103 1233 132 1330
rect 21 874 23 985
rect 23 874 49 985
rect 21 872 49 874
rect 261 1234 287 1332
rect 287 1234 290 1332
rect 175 873 202 987
rect 202 873 203 987
rect 416 1231 445 1331
rect 334 873 361 987
rect 361 873 362 987
rect 570 1231 604 1336
rect 495 873 522 987
rect 522 873 523 987
rect 727 1231 761 1334
rect 652 871 681 988
rect 887 1234 918 1330
rect 807 871 834 988
rect 834 871 836 988
rect 1044 1232 1076 1328
rect 970 872 997 988
rect 997 872 998 988
rect 1128 871 1155 987
rect 1155 871 1156 987
rect 79 419 107 530
rect 0 73 28 177
rect 159 79 187 183
rect 242 420 268 527
rect 268 420 270 527
rect 396 419 424 532
rect 319 73 347 184
rect 558 419 585 523
rect 585 419 587 523
rect 476 69 504 182
rect 715 419 741 520
rect 741 419 744 520
rect 634 184 664 185
rect 634 69 660 184
rect 660 69 664 184
rect 874 419 900 521
rect 900 419 902 521
rect 794 70 820 186
rect 820 70 822 186
rect 1030 419 1056 521
rect 1056 419 1058 521
rect 949 185 978 186
rect 949 71 976 185
rect 976 71 978 185
rect 1111 70 1137 187
rect 1137 70 1139 187
rect 1190 419 1216 521
rect 1216 419 1218 521
rect 1344 419 1372 525
rect 1270 70 1298 186
rect 1505 418 1533 525
rect 1425 68 1454 186
<< metal3 >>
rect 6 1336 1193 1352
rect 6 1332 570 1336
rect 6 1330 261 1332
rect 6 1233 103 1330
rect 132 1234 261 1330
rect 290 1331 570 1332
rect 290 1234 416 1331
rect 132 1233 416 1234
rect 6 1231 416 1233
rect 445 1231 570 1331
rect 604 1334 1193 1336
rect 604 1231 727 1334
rect 761 1330 1193 1334
rect 761 1234 887 1330
rect 918 1328 1193 1330
rect 918 1234 1044 1328
rect 761 1232 1044 1234
rect 1076 1232 1193 1328
rect 761 1231 1193 1232
rect 6 1226 1193 1231
rect 6 988 1193 992
rect 6 987 652 988
rect 6 985 175 987
rect 6 872 21 985
rect 49 873 175 985
rect 203 873 334 987
rect 362 873 495 987
rect 523 873 652 987
rect 49 872 652 873
rect 6 871 652 872
rect 681 871 807 988
rect 836 872 970 988
rect 998 987 1193 988
rect 998 872 1128 987
rect 836 871 1128 872
rect 1156 871 1193 987
rect 6 866 1193 871
rect -7 533 1534 541
rect -7 532 1537 533
rect -7 530 396 532
rect -7 419 79 530
rect 107 527 396 530
rect 107 420 242 527
rect 270 420 396 527
rect 107 419 396 420
rect 424 525 1537 532
rect 424 523 1344 525
rect 424 419 558 523
rect 587 521 1344 523
rect 587 520 874 521
rect 587 419 715 520
rect 744 419 874 520
rect 902 419 1030 521
rect 1058 419 1190 521
rect 1218 419 1344 521
rect 1372 419 1505 525
rect -7 418 1505 419
rect 1533 418 1537 525
rect -7 414 1537 418
rect 1501 413 1537 414
rect 1422 191 1458 192
rect -9 187 1532 191
rect -9 186 1111 187
rect -9 185 794 186
rect -9 184 634 185
rect -9 183 319 184
rect -9 177 159 183
rect -9 73 0 177
rect 28 79 159 177
rect 187 79 319 183
rect 28 73 319 79
rect 347 182 634 184
rect 347 73 476 182
rect -9 69 476 73
rect 504 69 634 182
rect 664 70 794 185
rect 822 71 949 186
rect 978 71 1111 186
rect 822 70 1111 71
rect 1139 186 1532 187
rect 1139 70 1270 186
rect 1298 70 1425 186
rect 664 69 1425 70
rect -9 68 1425 69
rect 1454 68 1532 186
rect -9 64 1532 68
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_0
timestamp 1717178954
transform 1 0 212 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_1
timestamp 1717178954
transform 1 0 54 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_2
timestamp 1717178954
transform 1 0 133 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_3
timestamp 1717178954
transform 1 0 449 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_4
timestamp 1717178954
transform 1 0 291 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_5
timestamp 1717178954
transform 1 0 370 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_6
timestamp 1717178954
transform 1 0 686 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_7
timestamp 1717178954
transform 1 0 528 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_8
timestamp 1717178954
transform 1 0 607 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_9
timestamp 1717178954
transform 1 0 923 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_10
timestamp 1717178954
transform 1 0 765 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_11
timestamp 1717178954
transform 1 0 844 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_12
timestamp 1717178954
transform 1 0 1081 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_13
timestamp 1717178954
transform 1 0 1002 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_14
timestamp 1717178954
transform 1 0 1476 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_15
timestamp 1717178954
transform 1 0 1160 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_16
timestamp 1717178954
transform 1 0 1239 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_17
timestamp 1717178954
transform 1 0 1318 0 1 294
box -54 -294 54 294
use sky130_fd_pr__nfet_01v8_U9XYXH  sky130_fd_pr__nfet_01v8_U9XYXH_18
timestamp 1717178954
transform 1 0 1397 0 1 294
box -54 -294 54 294
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_0
timestamp 1717178954
transform 1 0 72 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_1
timestamp 1717178954
transform 1 0 151 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_2
timestamp 1717178954
transform 1 0 230 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_3
timestamp 1717178954
transform 1 0 309 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_4
timestamp 1717178954
transform 1 0 388 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_5
timestamp 1717178954
transform 1 0 467 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_6
timestamp 1717178954
transform 1 0 546 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_7
timestamp 1717178954
transform 1 0 625 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_8
timestamp 1717178954
transform 1 0 704 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_9
timestamp 1717178954
transform 1 0 783 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_10
timestamp 1717178954
transform 1 0 862 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_11
timestamp 1717178954
transform 1 0 941 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_12
timestamp 1717178954
transform 1 0 1020 0 1 1100
box -72 -300 72 300
use sky130_fd_pr__pfet_01v8_lvt_YS6JVD  sky130_fd_pr__pfet_01v8_lvt_YS6JVD_13
timestamp 1717178954
transform 1 0 1099 0 1 1100
box -72 -300 72 300
<< labels >>
flabel metal1 -68 -63 70 -21 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 190 1413 300 1455 0 FreeSans 400 0 0 0 VCC
port 6 nsew
flabel metal3 1156 866 1193 992 0 FreeSans 400 0 0 0 OUT
port 7 nsew
flabel metal1 25 562 120 645 0 FreeSans 400 0 0 0 IBIAS
port 8 nsew
flabel metal1 43 738 138 834 0 FreeSans 400 0 0 0 DIFF_OUT
port 9 nsew
<< end >>
