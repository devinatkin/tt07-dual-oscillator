magic
tech sky130A
timestamp 1716419327
<< pwell >>
rect -834 -4855 834 4855
<< nmos >>
rect -736 -4750 -686 4750
rect -657 -4750 -607 4750
rect -578 -4750 -528 4750
rect -499 -4750 -449 4750
rect -420 -4750 -370 4750
rect -341 -4750 -291 4750
rect -262 -4750 -212 4750
rect -183 -4750 -133 4750
rect -104 -4750 -54 4750
rect -25 -4750 25 4750
rect 54 -4750 104 4750
rect 133 -4750 183 4750
rect 212 -4750 262 4750
rect 291 -4750 341 4750
rect 370 -4750 420 4750
rect 449 -4750 499 4750
rect 528 -4750 578 4750
rect 607 -4750 657 4750
rect 686 -4750 736 4750
<< ndiff >>
rect -765 4744 -736 4750
rect -765 -4744 -759 4744
rect -742 -4744 -736 4744
rect -765 -4750 -736 -4744
rect -686 4744 -657 4750
rect -686 -4744 -680 4744
rect -663 -4744 -657 4744
rect -686 -4750 -657 -4744
rect -607 4744 -578 4750
rect -607 -4744 -601 4744
rect -584 -4744 -578 4744
rect -607 -4750 -578 -4744
rect -528 4744 -499 4750
rect -528 -4744 -522 4744
rect -505 -4744 -499 4744
rect -528 -4750 -499 -4744
rect -449 4744 -420 4750
rect -449 -4744 -443 4744
rect -426 -4744 -420 4744
rect -449 -4750 -420 -4744
rect -370 4744 -341 4750
rect -370 -4744 -364 4744
rect -347 -4744 -341 4744
rect -370 -4750 -341 -4744
rect -291 4744 -262 4750
rect -291 -4744 -285 4744
rect -268 -4744 -262 4744
rect -291 -4750 -262 -4744
rect -212 4744 -183 4750
rect -212 -4744 -206 4744
rect -189 -4744 -183 4744
rect -212 -4750 -183 -4744
rect -133 4744 -104 4750
rect -133 -4744 -127 4744
rect -110 -4744 -104 4744
rect -133 -4750 -104 -4744
rect -54 4744 -25 4750
rect -54 -4744 -48 4744
rect -31 -4744 -25 4744
rect -54 -4750 -25 -4744
rect 25 4744 54 4750
rect 25 -4744 31 4744
rect 48 -4744 54 4744
rect 25 -4750 54 -4744
rect 104 4744 133 4750
rect 104 -4744 110 4744
rect 127 -4744 133 4744
rect 104 -4750 133 -4744
rect 183 4744 212 4750
rect 183 -4744 189 4744
rect 206 -4744 212 4744
rect 183 -4750 212 -4744
rect 262 4744 291 4750
rect 262 -4744 268 4744
rect 285 -4744 291 4744
rect 262 -4750 291 -4744
rect 341 4744 370 4750
rect 341 -4744 347 4744
rect 364 -4744 370 4744
rect 341 -4750 370 -4744
rect 420 4744 449 4750
rect 420 -4744 426 4744
rect 443 -4744 449 4744
rect 420 -4750 449 -4744
rect 499 4744 528 4750
rect 499 -4744 505 4744
rect 522 -4744 528 4744
rect 499 -4750 528 -4744
rect 578 4744 607 4750
rect 578 -4744 584 4744
rect 601 -4744 607 4744
rect 578 -4750 607 -4744
rect 657 4744 686 4750
rect 657 -4744 663 4744
rect 680 -4744 686 4744
rect 657 -4750 686 -4744
rect 736 4744 765 4750
rect 736 -4744 742 4744
rect 759 -4744 765 4744
rect 736 -4750 765 -4744
<< ndiffc >>
rect -759 -4744 -742 4744
rect -680 -4744 -663 4744
rect -601 -4744 -584 4744
rect -522 -4744 -505 4744
rect -443 -4744 -426 4744
rect -364 -4744 -347 4744
rect -285 -4744 -268 4744
rect -206 -4744 -189 4744
rect -127 -4744 -110 4744
rect -48 -4744 -31 4744
rect 31 -4744 48 4744
rect 110 -4744 127 4744
rect 189 -4744 206 4744
rect 268 -4744 285 4744
rect 347 -4744 364 4744
rect 426 -4744 443 4744
rect 505 -4744 522 4744
rect 584 -4744 601 4744
rect 663 -4744 680 4744
rect 742 -4744 759 4744
<< psubdiff >>
rect -816 4820 -768 4837
rect 768 4820 816 4837
rect -816 4789 -799 4820
rect 799 4789 816 4820
rect -816 -4820 -799 -4789
rect 799 -4820 816 -4789
rect -816 -4837 -768 -4820
rect 768 -4837 816 -4820
<< psubdiffcont >>
rect -768 4820 768 4837
rect -816 -4789 -799 4789
rect 799 -4789 816 4789
rect -768 -4837 768 -4820
<< poly >>
rect -736 4786 -686 4794
rect -736 4769 -728 4786
rect -694 4769 -686 4786
rect -736 4750 -686 4769
rect -657 4786 -607 4794
rect -657 4769 -649 4786
rect -615 4769 -607 4786
rect -657 4750 -607 4769
rect -578 4786 -528 4794
rect -578 4769 -570 4786
rect -536 4769 -528 4786
rect -578 4750 -528 4769
rect -499 4786 -449 4794
rect -499 4769 -491 4786
rect -457 4769 -449 4786
rect -499 4750 -449 4769
rect -420 4786 -370 4794
rect -420 4769 -412 4786
rect -378 4769 -370 4786
rect -420 4750 -370 4769
rect -341 4786 -291 4794
rect -341 4769 -333 4786
rect -299 4769 -291 4786
rect -341 4750 -291 4769
rect -262 4786 -212 4794
rect -262 4769 -254 4786
rect -220 4769 -212 4786
rect -262 4750 -212 4769
rect -183 4786 -133 4794
rect -183 4769 -175 4786
rect -141 4769 -133 4786
rect -183 4750 -133 4769
rect -104 4786 -54 4794
rect -104 4769 -96 4786
rect -62 4769 -54 4786
rect -104 4750 -54 4769
rect -25 4786 25 4794
rect -25 4769 -17 4786
rect 17 4769 25 4786
rect -25 4750 25 4769
rect 54 4786 104 4794
rect 54 4769 62 4786
rect 96 4769 104 4786
rect 54 4750 104 4769
rect 133 4786 183 4794
rect 133 4769 141 4786
rect 175 4769 183 4786
rect 133 4750 183 4769
rect 212 4786 262 4794
rect 212 4769 220 4786
rect 254 4769 262 4786
rect 212 4750 262 4769
rect 291 4786 341 4794
rect 291 4769 299 4786
rect 333 4769 341 4786
rect 291 4750 341 4769
rect 370 4786 420 4794
rect 370 4769 378 4786
rect 412 4769 420 4786
rect 370 4750 420 4769
rect 449 4786 499 4794
rect 449 4769 457 4786
rect 491 4769 499 4786
rect 449 4750 499 4769
rect 528 4786 578 4794
rect 528 4769 536 4786
rect 570 4769 578 4786
rect 528 4750 578 4769
rect 607 4786 657 4794
rect 607 4769 615 4786
rect 649 4769 657 4786
rect 607 4750 657 4769
rect 686 4786 736 4794
rect 686 4769 694 4786
rect 728 4769 736 4786
rect 686 4750 736 4769
rect -736 -4769 -686 -4750
rect -736 -4786 -728 -4769
rect -694 -4786 -686 -4769
rect -736 -4794 -686 -4786
rect -657 -4769 -607 -4750
rect -657 -4786 -649 -4769
rect -615 -4786 -607 -4769
rect -657 -4794 -607 -4786
rect -578 -4769 -528 -4750
rect -578 -4786 -570 -4769
rect -536 -4786 -528 -4769
rect -578 -4794 -528 -4786
rect -499 -4769 -449 -4750
rect -499 -4786 -491 -4769
rect -457 -4786 -449 -4769
rect -499 -4794 -449 -4786
rect -420 -4769 -370 -4750
rect -420 -4786 -412 -4769
rect -378 -4786 -370 -4769
rect -420 -4794 -370 -4786
rect -341 -4769 -291 -4750
rect -341 -4786 -333 -4769
rect -299 -4786 -291 -4769
rect -341 -4794 -291 -4786
rect -262 -4769 -212 -4750
rect -262 -4786 -254 -4769
rect -220 -4786 -212 -4769
rect -262 -4794 -212 -4786
rect -183 -4769 -133 -4750
rect -183 -4786 -175 -4769
rect -141 -4786 -133 -4769
rect -183 -4794 -133 -4786
rect -104 -4769 -54 -4750
rect -104 -4786 -96 -4769
rect -62 -4786 -54 -4769
rect -104 -4794 -54 -4786
rect -25 -4769 25 -4750
rect -25 -4786 -17 -4769
rect 17 -4786 25 -4769
rect -25 -4794 25 -4786
rect 54 -4769 104 -4750
rect 54 -4786 62 -4769
rect 96 -4786 104 -4769
rect 54 -4794 104 -4786
rect 133 -4769 183 -4750
rect 133 -4786 141 -4769
rect 175 -4786 183 -4769
rect 133 -4794 183 -4786
rect 212 -4769 262 -4750
rect 212 -4786 220 -4769
rect 254 -4786 262 -4769
rect 212 -4794 262 -4786
rect 291 -4769 341 -4750
rect 291 -4786 299 -4769
rect 333 -4786 341 -4769
rect 291 -4794 341 -4786
rect 370 -4769 420 -4750
rect 370 -4786 378 -4769
rect 412 -4786 420 -4769
rect 370 -4794 420 -4786
rect 449 -4769 499 -4750
rect 449 -4786 457 -4769
rect 491 -4786 499 -4769
rect 449 -4794 499 -4786
rect 528 -4769 578 -4750
rect 528 -4786 536 -4769
rect 570 -4786 578 -4769
rect 528 -4794 578 -4786
rect 607 -4769 657 -4750
rect 607 -4786 615 -4769
rect 649 -4786 657 -4769
rect 607 -4794 657 -4786
rect 686 -4769 736 -4750
rect 686 -4786 694 -4769
rect 728 -4786 736 -4769
rect 686 -4794 736 -4786
<< polycont >>
rect -728 4769 -694 4786
rect -649 4769 -615 4786
rect -570 4769 -536 4786
rect -491 4769 -457 4786
rect -412 4769 -378 4786
rect -333 4769 -299 4786
rect -254 4769 -220 4786
rect -175 4769 -141 4786
rect -96 4769 -62 4786
rect -17 4769 17 4786
rect 62 4769 96 4786
rect 141 4769 175 4786
rect 220 4769 254 4786
rect 299 4769 333 4786
rect 378 4769 412 4786
rect 457 4769 491 4786
rect 536 4769 570 4786
rect 615 4769 649 4786
rect 694 4769 728 4786
rect -728 -4786 -694 -4769
rect -649 -4786 -615 -4769
rect -570 -4786 -536 -4769
rect -491 -4786 -457 -4769
rect -412 -4786 -378 -4769
rect -333 -4786 -299 -4769
rect -254 -4786 -220 -4769
rect -175 -4786 -141 -4769
rect -96 -4786 -62 -4769
rect -17 -4786 17 -4769
rect 62 -4786 96 -4769
rect 141 -4786 175 -4769
rect 220 -4786 254 -4769
rect 299 -4786 333 -4769
rect 378 -4786 412 -4769
rect 457 -4786 491 -4769
rect 536 -4786 570 -4769
rect 615 -4786 649 -4769
rect 694 -4786 728 -4769
<< locali >>
rect -816 4820 -768 4837
rect 768 4820 816 4837
rect -816 4789 -799 4820
rect 799 4789 816 4820
rect -736 4769 -728 4786
rect -694 4769 -686 4786
rect -657 4769 -649 4786
rect -615 4769 -607 4786
rect -578 4769 -570 4786
rect -536 4769 -528 4786
rect -499 4769 -491 4786
rect -457 4769 -449 4786
rect -420 4769 -412 4786
rect -378 4769 -370 4786
rect -341 4769 -333 4786
rect -299 4769 -291 4786
rect -262 4769 -254 4786
rect -220 4769 -212 4786
rect -183 4769 -175 4786
rect -141 4769 -133 4786
rect -104 4769 -96 4786
rect -62 4769 -54 4786
rect -25 4769 -17 4786
rect 17 4769 25 4786
rect 54 4769 62 4786
rect 96 4769 104 4786
rect 133 4769 141 4786
rect 175 4769 183 4786
rect 212 4769 220 4786
rect 254 4769 262 4786
rect 291 4769 299 4786
rect 333 4769 341 4786
rect 370 4769 378 4786
rect 412 4769 420 4786
rect 449 4769 457 4786
rect 491 4769 499 4786
rect 528 4769 536 4786
rect 570 4769 578 4786
rect 607 4769 615 4786
rect 649 4769 657 4786
rect 686 4769 694 4786
rect 728 4769 736 4786
rect -759 4744 -742 4752
rect -759 -4752 -742 -4744
rect -680 4744 -663 4752
rect -680 -4752 -663 -4744
rect -601 4744 -584 4752
rect -601 -4752 -584 -4744
rect -522 4744 -505 4752
rect -522 -4752 -505 -4744
rect -443 4744 -426 4752
rect -443 -4752 -426 -4744
rect -364 4744 -347 4752
rect -364 -4752 -347 -4744
rect -285 4744 -268 4752
rect -285 -4752 -268 -4744
rect -206 4744 -189 4752
rect -206 -4752 -189 -4744
rect -127 4744 -110 4752
rect -127 -4752 -110 -4744
rect -48 4744 -31 4752
rect -48 -4752 -31 -4744
rect 31 4744 48 4752
rect 31 -4752 48 -4744
rect 110 4744 127 4752
rect 110 -4752 127 -4744
rect 189 4744 206 4752
rect 189 -4752 206 -4744
rect 268 4744 285 4752
rect 268 -4752 285 -4744
rect 347 4744 364 4752
rect 347 -4752 364 -4744
rect 426 4744 443 4752
rect 426 -4752 443 -4744
rect 505 4744 522 4752
rect 505 -4752 522 -4744
rect 584 4744 601 4752
rect 584 -4752 601 -4744
rect 663 4744 680 4752
rect 663 -4752 680 -4744
rect 742 4744 759 4752
rect 742 -4752 759 -4744
rect -736 -4786 -728 -4769
rect -694 -4786 -686 -4769
rect -657 -4786 -649 -4769
rect -615 -4786 -607 -4769
rect -578 -4786 -570 -4769
rect -536 -4786 -528 -4769
rect -499 -4786 -491 -4769
rect -457 -4786 -449 -4769
rect -420 -4786 -412 -4769
rect -378 -4786 -370 -4769
rect -341 -4786 -333 -4769
rect -299 -4786 -291 -4769
rect -262 -4786 -254 -4769
rect -220 -4786 -212 -4769
rect -183 -4786 -175 -4769
rect -141 -4786 -133 -4769
rect -104 -4786 -96 -4769
rect -62 -4786 -54 -4769
rect -25 -4786 -17 -4769
rect 17 -4786 25 -4769
rect 54 -4786 62 -4769
rect 96 -4786 104 -4769
rect 133 -4786 141 -4769
rect 175 -4786 183 -4769
rect 212 -4786 220 -4769
rect 254 -4786 262 -4769
rect 291 -4786 299 -4769
rect 333 -4786 341 -4769
rect 370 -4786 378 -4769
rect 412 -4786 420 -4769
rect 449 -4786 457 -4769
rect 491 -4786 499 -4769
rect 528 -4786 536 -4769
rect 570 -4786 578 -4769
rect 607 -4786 615 -4769
rect 649 -4786 657 -4769
rect 686 -4786 694 -4769
rect 728 -4786 736 -4769
rect -816 -4820 -799 -4789
rect 799 -4820 816 -4789
rect -816 -4837 -768 -4820
rect 768 -4837 816 -4820
<< viali >>
rect -728 4769 -694 4786
rect -649 4769 -615 4786
rect -570 4769 -536 4786
rect -491 4769 -457 4786
rect -412 4769 -378 4786
rect -333 4769 -299 4786
rect -254 4769 -220 4786
rect -175 4769 -141 4786
rect -96 4769 -62 4786
rect -17 4769 17 4786
rect 62 4769 96 4786
rect 141 4769 175 4786
rect 220 4769 254 4786
rect 299 4769 333 4786
rect 378 4769 412 4786
rect 457 4769 491 4786
rect 536 4769 570 4786
rect 615 4769 649 4786
rect 694 4769 728 4786
rect -759 -4744 -742 4744
rect -680 -4744 -663 4744
rect -601 -4744 -584 4744
rect -522 -4744 -505 4744
rect -443 -4744 -426 4744
rect -364 -4744 -347 4744
rect -285 -4744 -268 4744
rect -206 -4744 -189 4744
rect -127 -4744 -110 4744
rect -48 -4744 -31 4744
rect 31 -4744 48 4744
rect 110 -4744 127 4744
rect 189 -4744 206 4744
rect 268 -4744 285 4744
rect 347 -4744 364 4744
rect 426 -4744 443 4744
rect 505 -4744 522 4744
rect 584 -4744 601 4744
rect 663 -4744 680 4744
rect 742 -4744 759 4744
rect -728 -4786 -694 -4769
rect -649 -4786 -615 -4769
rect -570 -4786 -536 -4769
rect -491 -4786 -457 -4769
rect -412 -4786 -378 -4769
rect -333 -4786 -299 -4769
rect -254 -4786 -220 -4769
rect -175 -4786 -141 -4769
rect -96 -4786 -62 -4769
rect -17 -4786 17 -4769
rect 62 -4786 96 -4769
rect 141 -4786 175 -4769
rect 220 -4786 254 -4769
rect 299 -4786 333 -4769
rect 378 -4786 412 -4769
rect 457 -4786 491 -4769
rect 536 -4786 570 -4769
rect 615 -4786 649 -4769
rect 694 -4786 728 -4769
<< metal1 >>
rect -734 4786 -688 4789
rect -734 4769 -728 4786
rect -694 4769 -688 4786
rect -734 4766 -688 4769
rect -655 4786 -609 4789
rect -655 4769 -649 4786
rect -615 4769 -609 4786
rect -655 4766 -609 4769
rect -576 4786 -530 4789
rect -576 4769 -570 4786
rect -536 4769 -530 4786
rect -576 4766 -530 4769
rect -497 4786 -451 4789
rect -497 4769 -491 4786
rect -457 4769 -451 4786
rect -497 4766 -451 4769
rect -418 4786 -372 4789
rect -418 4769 -412 4786
rect -378 4769 -372 4786
rect -418 4766 -372 4769
rect -339 4786 -293 4789
rect -339 4769 -333 4786
rect -299 4769 -293 4786
rect -339 4766 -293 4769
rect -260 4786 -214 4789
rect -260 4769 -254 4786
rect -220 4769 -214 4786
rect -260 4766 -214 4769
rect -181 4786 -135 4789
rect -181 4769 -175 4786
rect -141 4769 -135 4786
rect -181 4766 -135 4769
rect -102 4786 -56 4789
rect -102 4769 -96 4786
rect -62 4769 -56 4786
rect -102 4766 -56 4769
rect -23 4786 23 4789
rect -23 4769 -17 4786
rect 17 4769 23 4786
rect -23 4766 23 4769
rect 56 4786 102 4789
rect 56 4769 62 4786
rect 96 4769 102 4786
rect 56 4766 102 4769
rect 135 4786 181 4789
rect 135 4769 141 4786
rect 175 4769 181 4786
rect 135 4766 181 4769
rect 214 4786 260 4789
rect 214 4769 220 4786
rect 254 4769 260 4786
rect 214 4766 260 4769
rect 293 4786 339 4789
rect 293 4769 299 4786
rect 333 4769 339 4786
rect 293 4766 339 4769
rect 372 4786 418 4789
rect 372 4769 378 4786
rect 412 4769 418 4786
rect 372 4766 418 4769
rect 451 4786 497 4789
rect 451 4769 457 4786
rect 491 4769 497 4786
rect 451 4766 497 4769
rect 530 4786 576 4789
rect 530 4769 536 4786
rect 570 4769 576 4786
rect 530 4766 576 4769
rect 609 4786 655 4789
rect 609 4769 615 4786
rect 649 4769 655 4786
rect 609 4766 655 4769
rect 688 4786 734 4789
rect 688 4769 694 4786
rect 728 4769 734 4786
rect 688 4766 734 4769
rect -762 4744 -739 4750
rect -762 -4744 -759 4744
rect -742 -4744 -739 4744
rect -762 -4750 -739 -4744
rect -683 4744 -660 4750
rect -683 -4744 -680 4744
rect -663 -4744 -660 4744
rect -683 -4750 -660 -4744
rect -604 4744 -581 4750
rect -604 -4744 -601 4744
rect -584 -4744 -581 4744
rect -604 -4750 -581 -4744
rect -525 4744 -502 4750
rect -525 -4744 -522 4744
rect -505 -4744 -502 4744
rect -525 -4750 -502 -4744
rect -446 4744 -423 4750
rect -446 -4744 -443 4744
rect -426 -4744 -423 4744
rect -446 -4750 -423 -4744
rect -367 4744 -344 4750
rect -367 -4744 -364 4744
rect -347 -4744 -344 4744
rect -367 -4750 -344 -4744
rect -288 4744 -265 4750
rect -288 -4744 -285 4744
rect -268 -4744 -265 4744
rect -288 -4750 -265 -4744
rect -209 4744 -186 4750
rect -209 -4744 -206 4744
rect -189 -4744 -186 4744
rect -209 -4750 -186 -4744
rect -130 4744 -107 4750
rect -130 -4744 -127 4744
rect -110 -4744 -107 4744
rect -130 -4750 -107 -4744
rect -51 4744 -28 4750
rect -51 -4744 -48 4744
rect -31 -4744 -28 4744
rect -51 -4750 -28 -4744
rect 28 4744 51 4750
rect 28 -4744 31 4744
rect 48 -4744 51 4744
rect 28 -4750 51 -4744
rect 107 4744 130 4750
rect 107 -4744 110 4744
rect 127 -4744 130 4744
rect 107 -4750 130 -4744
rect 186 4744 209 4750
rect 186 -4744 189 4744
rect 206 -4744 209 4744
rect 186 -4750 209 -4744
rect 265 4744 288 4750
rect 265 -4744 268 4744
rect 285 -4744 288 4744
rect 265 -4750 288 -4744
rect 344 4744 367 4750
rect 344 -4744 347 4744
rect 364 -4744 367 4744
rect 344 -4750 367 -4744
rect 423 4744 446 4750
rect 423 -4744 426 4744
rect 443 -4744 446 4744
rect 423 -4750 446 -4744
rect 502 4744 525 4750
rect 502 -4744 505 4744
rect 522 -4744 525 4744
rect 502 -4750 525 -4744
rect 581 4744 604 4750
rect 581 -4744 584 4744
rect 601 -4744 604 4744
rect 581 -4750 604 -4744
rect 660 4744 683 4750
rect 660 -4744 663 4744
rect 680 -4744 683 4744
rect 660 -4750 683 -4744
rect 739 4744 762 4750
rect 739 -4744 742 4744
rect 759 -4744 762 4744
rect 739 -4750 762 -4744
rect -734 -4769 -688 -4766
rect -734 -4786 -728 -4769
rect -694 -4786 -688 -4769
rect -734 -4789 -688 -4786
rect -655 -4769 -609 -4766
rect -655 -4786 -649 -4769
rect -615 -4786 -609 -4769
rect -655 -4789 -609 -4786
rect -576 -4769 -530 -4766
rect -576 -4786 -570 -4769
rect -536 -4786 -530 -4769
rect -576 -4789 -530 -4786
rect -497 -4769 -451 -4766
rect -497 -4786 -491 -4769
rect -457 -4786 -451 -4769
rect -497 -4789 -451 -4786
rect -418 -4769 -372 -4766
rect -418 -4786 -412 -4769
rect -378 -4786 -372 -4769
rect -418 -4789 -372 -4786
rect -339 -4769 -293 -4766
rect -339 -4786 -333 -4769
rect -299 -4786 -293 -4769
rect -339 -4789 -293 -4786
rect -260 -4769 -214 -4766
rect -260 -4786 -254 -4769
rect -220 -4786 -214 -4769
rect -260 -4789 -214 -4786
rect -181 -4769 -135 -4766
rect -181 -4786 -175 -4769
rect -141 -4786 -135 -4769
rect -181 -4789 -135 -4786
rect -102 -4769 -56 -4766
rect -102 -4786 -96 -4769
rect -62 -4786 -56 -4769
rect -102 -4789 -56 -4786
rect -23 -4769 23 -4766
rect -23 -4786 -17 -4769
rect 17 -4786 23 -4769
rect -23 -4789 23 -4786
rect 56 -4769 102 -4766
rect 56 -4786 62 -4769
rect 96 -4786 102 -4769
rect 56 -4789 102 -4786
rect 135 -4769 181 -4766
rect 135 -4786 141 -4769
rect 175 -4786 181 -4769
rect 135 -4789 181 -4786
rect 214 -4769 260 -4766
rect 214 -4786 220 -4769
rect 254 -4786 260 -4769
rect 214 -4789 260 -4786
rect 293 -4769 339 -4766
rect 293 -4786 299 -4769
rect 333 -4786 339 -4769
rect 293 -4789 339 -4786
rect 372 -4769 418 -4766
rect 372 -4786 378 -4769
rect 412 -4786 418 -4769
rect 372 -4789 418 -4786
rect 451 -4769 497 -4766
rect 451 -4786 457 -4769
rect 491 -4786 497 -4769
rect 451 -4789 497 -4786
rect 530 -4769 576 -4766
rect 530 -4786 536 -4769
rect 570 -4786 576 -4769
rect 530 -4789 576 -4786
rect 609 -4769 655 -4766
rect 609 -4786 615 -4769
rect 649 -4786 655 -4769
rect 609 -4789 655 -4786
rect 688 -4769 734 -4766
rect 688 -4786 694 -4769
rect 728 -4786 734 -4769
rect 688 -4789 734 -4786
<< properties >>
string FIXED_BBOX -807 -4828 807 4828
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 95.0 l 0.5 m 1 nf 19 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
