magic
tech sky130A
timestamp 1716325537
<< pwell >>
rect -123 -5836 123 5836
<< nmos >>
rect -25 5231 25 5731
rect -25 4622 25 5122
rect -25 4013 25 4513
rect -25 3404 25 3904
rect -25 2795 25 3295
rect -25 2186 25 2686
rect -25 1577 25 2077
rect -25 968 25 1468
rect -25 359 25 859
rect -25 -250 25 250
rect -25 -859 25 -359
rect -25 -1468 25 -968
rect -25 -2077 25 -1577
rect -25 -2686 25 -2186
rect -25 -3295 25 -2795
rect -25 -3904 25 -3404
rect -25 -4513 25 -4013
rect -25 -5122 25 -4622
rect -25 -5731 25 -5231
<< ndiff >>
rect -54 5725 -25 5731
rect -54 5237 -48 5725
rect -31 5237 -25 5725
rect -54 5231 -25 5237
rect 25 5725 54 5731
rect 25 5237 31 5725
rect 48 5237 54 5725
rect 25 5231 54 5237
rect -54 5116 -25 5122
rect -54 4628 -48 5116
rect -31 4628 -25 5116
rect -54 4622 -25 4628
rect 25 5116 54 5122
rect 25 4628 31 5116
rect 48 4628 54 5116
rect 25 4622 54 4628
rect -54 4507 -25 4513
rect -54 4019 -48 4507
rect -31 4019 -25 4507
rect -54 4013 -25 4019
rect 25 4507 54 4513
rect 25 4019 31 4507
rect 48 4019 54 4507
rect 25 4013 54 4019
rect -54 3898 -25 3904
rect -54 3410 -48 3898
rect -31 3410 -25 3898
rect -54 3404 -25 3410
rect 25 3898 54 3904
rect 25 3410 31 3898
rect 48 3410 54 3898
rect 25 3404 54 3410
rect -54 3289 -25 3295
rect -54 2801 -48 3289
rect -31 2801 -25 3289
rect -54 2795 -25 2801
rect 25 3289 54 3295
rect 25 2801 31 3289
rect 48 2801 54 3289
rect 25 2795 54 2801
rect -54 2680 -25 2686
rect -54 2192 -48 2680
rect -31 2192 -25 2680
rect -54 2186 -25 2192
rect 25 2680 54 2686
rect 25 2192 31 2680
rect 48 2192 54 2680
rect 25 2186 54 2192
rect -54 2071 -25 2077
rect -54 1583 -48 2071
rect -31 1583 -25 2071
rect -54 1577 -25 1583
rect 25 2071 54 2077
rect 25 1583 31 2071
rect 48 1583 54 2071
rect 25 1577 54 1583
rect -54 1462 -25 1468
rect -54 974 -48 1462
rect -31 974 -25 1462
rect -54 968 -25 974
rect 25 1462 54 1468
rect 25 974 31 1462
rect 48 974 54 1462
rect 25 968 54 974
rect -54 853 -25 859
rect -54 365 -48 853
rect -31 365 -25 853
rect -54 359 -25 365
rect 25 853 54 859
rect 25 365 31 853
rect 48 365 54 853
rect 25 359 54 365
rect -54 244 -25 250
rect -54 -244 -48 244
rect -31 -244 -25 244
rect -54 -250 -25 -244
rect 25 244 54 250
rect 25 -244 31 244
rect 48 -244 54 244
rect 25 -250 54 -244
rect -54 -365 -25 -359
rect -54 -853 -48 -365
rect -31 -853 -25 -365
rect -54 -859 -25 -853
rect 25 -365 54 -359
rect 25 -853 31 -365
rect 48 -853 54 -365
rect 25 -859 54 -853
rect -54 -974 -25 -968
rect -54 -1462 -48 -974
rect -31 -1462 -25 -974
rect -54 -1468 -25 -1462
rect 25 -974 54 -968
rect 25 -1462 31 -974
rect 48 -1462 54 -974
rect 25 -1468 54 -1462
rect -54 -1583 -25 -1577
rect -54 -2071 -48 -1583
rect -31 -2071 -25 -1583
rect -54 -2077 -25 -2071
rect 25 -1583 54 -1577
rect 25 -2071 31 -1583
rect 48 -2071 54 -1583
rect 25 -2077 54 -2071
rect -54 -2192 -25 -2186
rect -54 -2680 -48 -2192
rect -31 -2680 -25 -2192
rect -54 -2686 -25 -2680
rect 25 -2192 54 -2186
rect 25 -2680 31 -2192
rect 48 -2680 54 -2192
rect 25 -2686 54 -2680
rect -54 -2801 -25 -2795
rect -54 -3289 -48 -2801
rect -31 -3289 -25 -2801
rect -54 -3295 -25 -3289
rect 25 -2801 54 -2795
rect 25 -3289 31 -2801
rect 48 -3289 54 -2801
rect 25 -3295 54 -3289
rect -54 -3410 -25 -3404
rect -54 -3898 -48 -3410
rect -31 -3898 -25 -3410
rect -54 -3904 -25 -3898
rect 25 -3410 54 -3404
rect 25 -3898 31 -3410
rect 48 -3898 54 -3410
rect 25 -3904 54 -3898
rect -54 -4019 -25 -4013
rect -54 -4507 -48 -4019
rect -31 -4507 -25 -4019
rect -54 -4513 -25 -4507
rect 25 -4019 54 -4013
rect 25 -4507 31 -4019
rect 48 -4507 54 -4019
rect 25 -4513 54 -4507
rect -54 -4628 -25 -4622
rect -54 -5116 -48 -4628
rect -31 -5116 -25 -4628
rect -54 -5122 -25 -5116
rect 25 -4628 54 -4622
rect 25 -5116 31 -4628
rect 48 -5116 54 -4628
rect 25 -5122 54 -5116
rect -54 -5237 -25 -5231
rect -54 -5725 -48 -5237
rect -31 -5725 -25 -5237
rect -54 -5731 -25 -5725
rect 25 -5237 54 -5231
rect 25 -5725 31 -5237
rect 48 -5725 54 -5237
rect 25 -5731 54 -5725
<< ndiffc >>
rect -48 5237 -31 5725
rect 31 5237 48 5725
rect -48 4628 -31 5116
rect 31 4628 48 5116
rect -48 4019 -31 4507
rect 31 4019 48 4507
rect -48 3410 -31 3898
rect 31 3410 48 3898
rect -48 2801 -31 3289
rect 31 2801 48 3289
rect -48 2192 -31 2680
rect 31 2192 48 2680
rect -48 1583 -31 2071
rect 31 1583 48 2071
rect -48 974 -31 1462
rect 31 974 48 1462
rect -48 365 -31 853
rect 31 365 48 853
rect -48 -244 -31 244
rect 31 -244 48 244
rect -48 -853 -31 -365
rect 31 -853 48 -365
rect -48 -1462 -31 -974
rect 31 -1462 48 -974
rect -48 -2071 -31 -1583
rect 31 -2071 48 -1583
rect -48 -2680 -31 -2192
rect 31 -2680 48 -2192
rect -48 -3289 -31 -2801
rect 31 -3289 48 -2801
rect -48 -3898 -31 -3410
rect 31 -3898 48 -3410
rect -48 -4507 -31 -4019
rect 31 -4507 48 -4019
rect -48 -5116 -31 -4628
rect 31 -5116 48 -4628
rect -48 -5725 -31 -5237
rect 31 -5725 48 -5237
<< psubdiff >>
rect -105 5801 -57 5818
rect 57 5801 105 5818
rect -105 5770 -88 5801
rect 88 5770 105 5801
rect -105 -5801 -88 -5770
rect 88 -5801 105 -5770
rect -105 -5818 -57 -5801
rect 57 -5818 105 -5801
<< psubdiffcont >>
rect -57 5801 57 5818
rect -105 -5770 -88 5770
rect 88 -5770 105 5770
rect -57 -5818 57 -5801
<< poly >>
rect -25 5767 25 5775
rect -25 5750 -17 5767
rect 17 5750 25 5767
rect -25 5731 25 5750
rect -25 5212 25 5231
rect -25 5195 -17 5212
rect 17 5195 25 5212
rect -25 5187 25 5195
rect -25 5158 25 5166
rect -25 5141 -17 5158
rect 17 5141 25 5158
rect -25 5122 25 5141
rect -25 4603 25 4622
rect -25 4586 -17 4603
rect 17 4586 25 4603
rect -25 4578 25 4586
rect -25 4549 25 4557
rect -25 4532 -17 4549
rect 17 4532 25 4549
rect -25 4513 25 4532
rect -25 3994 25 4013
rect -25 3977 -17 3994
rect 17 3977 25 3994
rect -25 3969 25 3977
rect -25 3940 25 3948
rect -25 3923 -17 3940
rect 17 3923 25 3940
rect -25 3904 25 3923
rect -25 3385 25 3404
rect -25 3368 -17 3385
rect 17 3368 25 3385
rect -25 3360 25 3368
rect -25 3331 25 3339
rect -25 3314 -17 3331
rect 17 3314 25 3331
rect -25 3295 25 3314
rect -25 2776 25 2795
rect -25 2759 -17 2776
rect 17 2759 25 2776
rect -25 2751 25 2759
rect -25 2722 25 2730
rect -25 2705 -17 2722
rect 17 2705 25 2722
rect -25 2686 25 2705
rect -25 2167 25 2186
rect -25 2150 -17 2167
rect 17 2150 25 2167
rect -25 2142 25 2150
rect -25 2113 25 2121
rect -25 2096 -17 2113
rect 17 2096 25 2113
rect -25 2077 25 2096
rect -25 1558 25 1577
rect -25 1541 -17 1558
rect 17 1541 25 1558
rect -25 1533 25 1541
rect -25 1504 25 1512
rect -25 1487 -17 1504
rect 17 1487 25 1504
rect -25 1468 25 1487
rect -25 949 25 968
rect -25 932 -17 949
rect 17 932 25 949
rect -25 924 25 932
rect -25 895 25 903
rect -25 878 -17 895
rect 17 878 25 895
rect -25 859 25 878
rect -25 340 25 359
rect -25 323 -17 340
rect 17 323 25 340
rect -25 315 25 323
rect -25 286 25 294
rect -25 269 -17 286
rect 17 269 25 286
rect -25 250 25 269
rect -25 -269 25 -250
rect -25 -286 -17 -269
rect 17 -286 25 -269
rect -25 -294 25 -286
rect -25 -323 25 -315
rect -25 -340 -17 -323
rect 17 -340 25 -323
rect -25 -359 25 -340
rect -25 -878 25 -859
rect -25 -895 -17 -878
rect 17 -895 25 -878
rect -25 -903 25 -895
rect -25 -932 25 -924
rect -25 -949 -17 -932
rect 17 -949 25 -932
rect -25 -968 25 -949
rect -25 -1487 25 -1468
rect -25 -1504 -17 -1487
rect 17 -1504 25 -1487
rect -25 -1512 25 -1504
rect -25 -1541 25 -1533
rect -25 -1558 -17 -1541
rect 17 -1558 25 -1541
rect -25 -1577 25 -1558
rect -25 -2096 25 -2077
rect -25 -2113 -17 -2096
rect 17 -2113 25 -2096
rect -25 -2121 25 -2113
rect -25 -2150 25 -2142
rect -25 -2167 -17 -2150
rect 17 -2167 25 -2150
rect -25 -2186 25 -2167
rect -25 -2705 25 -2686
rect -25 -2722 -17 -2705
rect 17 -2722 25 -2705
rect -25 -2730 25 -2722
rect -25 -2759 25 -2751
rect -25 -2776 -17 -2759
rect 17 -2776 25 -2759
rect -25 -2795 25 -2776
rect -25 -3314 25 -3295
rect -25 -3331 -17 -3314
rect 17 -3331 25 -3314
rect -25 -3339 25 -3331
rect -25 -3368 25 -3360
rect -25 -3385 -17 -3368
rect 17 -3385 25 -3368
rect -25 -3404 25 -3385
rect -25 -3923 25 -3904
rect -25 -3940 -17 -3923
rect 17 -3940 25 -3923
rect -25 -3948 25 -3940
rect -25 -3977 25 -3969
rect -25 -3994 -17 -3977
rect 17 -3994 25 -3977
rect -25 -4013 25 -3994
rect -25 -4532 25 -4513
rect -25 -4549 -17 -4532
rect 17 -4549 25 -4532
rect -25 -4557 25 -4549
rect -25 -4586 25 -4578
rect -25 -4603 -17 -4586
rect 17 -4603 25 -4586
rect -25 -4622 25 -4603
rect -25 -5141 25 -5122
rect -25 -5158 -17 -5141
rect 17 -5158 25 -5141
rect -25 -5166 25 -5158
rect -25 -5195 25 -5187
rect -25 -5212 -17 -5195
rect 17 -5212 25 -5195
rect -25 -5231 25 -5212
rect -25 -5750 25 -5731
rect -25 -5767 -17 -5750
rect 17 -5767 25 -5750
rect -25 -5775 25 -5767
<< polycont >>
rect -17 5750 17 5767
rect -17 5195 17 5212
rect -17 5141 17 5158
rect -17 4586 17 4603
rect -17 4532 17 4549
rect -17 3977 17 3994
rect -17 3923 17 3940
rect -17 3368 17 3385
rect -17 3314 17 3331
rect -17 2759 17 2776
rect -17 2705 17 2722
rect -17 2150 17 2167
rect -17 2096 17 2113
rect -17 1541 17 1558
rect -17 1487 17 1504
rect -17 932 17 949
rect -17 878 17 895
rect -17 323 17 340
rect -17 269 17 286
rect -17 -286 17 -269
rect -17 -340 17 -323
rect -17 -895 17 -878
rect -17 -949 17 -932
rect -17 -1504 17 -1487
rect -17 -1558 17 -1541
rect -17 -2113 17 -2096
rect -17 -2167 17 -2150
rect -17 -2722 17 -2705
rect -17 -2776 17 -2759
rect -17 -3331 17 -3314
rect -17 -3385 17 -3368
rect -17 -3940 17 -3923
rect -17 -3994 17 -3977
rect -17 -4549 17 -4532
rect -17 -4603 17 -4586
rect -17 -5158 17 -5141
rect -17 -5212 17 -5195
rect -17 -5767 17 -5750
<< locali >>
rect -105 5801 -57 5818
rect 57 5801 105 5818
rect -105 5770 -88 5801
rect 88 5770 105 5801
rect -25 5750 -17 5767
rect 17 5750 25 5767
rect -48 5725 -31 5733
rect -48 5229 -31 5237
rect 31 5725 48 5733
rect 31 5229 48 5237
rect -25 5195 -17 5212
rect 17 5195 25 5212
rect -25 5141 -17 5158
rect 17 5141 25 5158
rect -48 5116 -31 5124
rect -48 4620 -31 4628
rect 31 5116 48 5124
rect 31 4620 48 4628
rect -25 4586 -17 4603
rect 17 4586 25 4603
rect -25 4532 -17 4549
rect 17 4532 25 4549
rect -48 4507 -31 4515
rect -48 4011 -31 4019
rect 31 4507 48 4515
rect 31 4011 48 4019
rect -25 3977 -17 3994
rect 17 3977 25 3994
rect -25 3923 -17 3940
rect 17 3923 25 3940
rect -48 3898 -31 3906
rect -48 3402 -31 3410
rect 31 3898 48 3906
rect 31 3402 48 3410
rect -25 3368 -17 3385
rect 17 3368 25 3385
rect -25 3314 -17 3331
rect 17 3314 25 3331
rect -48 3289 -31 3297
rect -48 2793 -31 2801
rect 31 3289 48 3297
rect 31 2793 48 2801
rect -25 2759 -17 2776
rect 17 2759 25 2776
rect -25 2705 -17 2722
rect 17 2705 25 2722
rect -48 2680 -31 2688
rect -48 2184 -31 2192
rect 31 2680 48 2688
rect 31 2184 48 2192
rect -25 2150 -17 2167
rect 17 2150 25 2167
rect -25 2096 -17 2113
rect 17 2096 25 2113
rect -48 2071 -31 2079
rect -48 1575 -31 1583
rect 31 2071 48 2079
rect 31 1575 48 1583
rect -25 1541 -17 1558
rect 17 1541 25 1558
rect -25 1487 -17 1504
rect 17 1487 25 1504
rect -48 1462 -31 1470
rect -48 966 -31 974
rect 31 1462 48 1470
rect 31 966 48 974
rect -25 932 -17 949
rect 17 932 25 949
rect -25 878 -17 895
rect 17 878 25 895
rect -48 853 -31 861
rect -48 357 -31 365
rect 31 853 48 861
rect 31 357 48 365
rect -25 323 -17 340
rect 17 323 25 340
rect -25 269 -17 286
rect 17 269 25 286
rect -48 244 -31 252
rect -48 -252 -31 -244
rect 31 244 48 252
rect 31 -252 48 -244
rect -25 -286 -17 -269
rect 17 -286 25 -269
rect -25 -340 -17 -323
rect 17 -340 25 -323
rect -48 -365 -31 -357
rect -48 -861 -31 -853
rect 31 -365 48 -357
rect 31 -861 48 -853
rect -25 -895 -17 -878
rect 17 -895 25 -878
rect -25 -949 -17 -932
rect 17 -949 25 -932
rect -48 -974 -31 -966
rect -48 -1470 -31 -1462
rect 31 -974 48 -966
rect 31 -1470 48 -1462
rect -25 -1504 -17 -1487
rect 17 -1504 25 -1487
rect -25 -1558 -17 -1541
rect 17 -1558 25 -1541
rect -48 -1583 -31 -1575
rect -48 -2079 -31 -2071
rect 31 -1583 48 -1575
rect 31 -2079 48 -2071
rect -25 -2113 -17 -2096
rect 17 -2113 25 -2096
rect -25 -2167 -17 -2150
rect 17 -2167 25 -2150
rect -48 -2192 -31 -2184
rect -48 -2688 -31 -2680
rect 31 -2192 48 -2184
rect 31 -2688 48 -2680
rect -25 -2722 -17 -2705
rect 17 -2722 25 -2705
rect -25 -2776 -17 -2759
rect 17 -2776 25 -2759
rect -48 -2801 -31 -2793
rect -48 -3297 -31 -3289
rect 31 -2801 48 -2793
rect 31 -3297 48 -3289
rect -25 -3331 -17 -3314
rect 17 -3331 25 -3314
rect -25 -3385 -17 -3368
rect 17 -3385 25 -3368
rect -48 -3410 -31 -3402
rect -48 -3906 -31 -3898
rect 31 -3410 48 -3402
rect 31 -3906 48 -3898
rect -25 -3940 -17 -3923
rect 17 -3940 25 -3923
rect -25 -3994 -17 -3977
rect 17 -3994 25 -3977
rect -48 -4019 -31 -4011
rect -48 -4515 -31 -4507
rect 31 -4019 48 -4011
rect 31 -4515 48 -4507
rect -25 -4549 -17 -4532
rect 17 -4549 25 -4532
rect -25 -4603 -17 -4586
rect 17 -4603 25 -4586
rect -48 -4628 -31 -4620
rect -48 -5124 -31 -5116
rect 31 -4628 48 -4620
rect 31 -5124 48 -5116
rect -25 -5158 -17 -5141
rect 17 -5158 25 -5141
rect -25 -5212 -17 -5195
rect 17 -5212 25 -5195
rect -48 -5237 -31 -5229
rect -48 -5733 -31 -5725
rect 31 -5237 48 -5229
rect 31 -5733 48 -5725
rect -25 -5767 -17 -5750
rect 17 -5767 25 -5750
rect -105 -5801 -88 -5770
rect 88 -5801 105 -5770
rect -105 -5818 -57 -5801
rect 57 -5818 105 -5801
<< viali >>
rect -17 5750 17 5767
rect -48 5237 -31 5725
rect 31 5237 48 5725
rect -17 5195 17 5212
rect -17 5141 17 5158
rect -48 4628 -31 5116
rect 31 4628 48 5116
rect -17 4586 17 4603
rect -17 4532 17 4549
rect -48 4019 -31 4507
rect 31 4019 48 4507
rect -17 3977 17 3994
rect -17 3923 17 3940
rect -48 3410 -31 3898
rect 31 3410 48 3898
rect -17 3368 17 3385
rect -17 3314 17 3331
rect -48 2801 -31 3289
rect 31 2801 48 3289
rect -17 2759 17 2776
rect -17 2705 17 2722
rect -48 2192 -31 2680
rect 31 2192 48 2680
rect -17 2150 17 2167
rect -17 2096 17 2113
rect -48 1583 -31 2071
rect 31 1583 48 2071
rect -17 1541 17 1558
rect -17 1487 17 1504
rect -48 974 -31 1462
rect 31 974 48 1462
rect -17 932 17 949
rect -17 878 17 895
rect -48 365 -31 853
rect 31 365 48 853
rect -17 323 17 340
rect -17 269 17 286
rect -48 -244 -31 244
rect 31 -244 48 244
rect -17 -286 17 -269
rect -17 -340 17 -323
rect -48 -853 -31 -365
rect 31 -853 48 -365
rect -17 -895 17 -878
rect -17 -949 17 -932
rect -48 -1462 -31 -974
rect 31 -1462 48 -974
rect -17 -1504 17 -1487
rect -17 -1558 17 -1541
rect -48 -2071 -31 -1583
rect 31 -2071 48 -1583
rect -17 -2113 17 -2096
rect -17 -2167 17 -2150
rect -48 -2680 -31 -2192
rect 31 -2680 48 -2192
rect -17 -2722 17 -2705
rect -17 -2776 17 -2759
rect -48 -3289 -31 -2801
rect 31 -3289 48 -2801
rect -17 -3331 17 -3314
rect -17 -3385 17 -3368
rect -48 -3898 -31 -3410
rect 31 -3898 48 -3410
rect -17 -3940 17 -3923
rect -17 -3994 17 -3977
rect -48 -4507 -31 -4019
rect 31 -4507 48 -4019
rect -17 -4549 17 -4532
rect -17 -4603 17 -4586
rect -48 -5116 -31 -4628
rect 31 -5116 48 -4628
rect -17 -5158 17 -5141
rect -17 -5212 17 -5195
rect -48 -5725 -31 -5237
rect 31 -5725 48 -5237
rect -17 -5767 17 -5750
<< metal1 >>
rect -23 5767 23 5770
rect -23 5750 -17 5767
rect 17 5750 23 5767
rect -23 5747 23 5750
rect -51 5725 -28 5731
rect -51 5237 -48 5725
rect -31 5237 -28 5725
rect -51 5231 -28 5237
rect 28 5725 51 5731
rect 28 5237 31 5725
rect 48 5237 51 5725
rect 28 5231 51 5237
rect -23 5212 23 5215
rect -23 5195 -17 5212
rect 17 5195 23 5212
rect -23 5192 23 5195
rect -23 5158 23 5161
rect -23 5141 -17 5158
rect 17 5141 23 5158
rect -23 5138 23 5141
rect -51 5116 -28 5122
rect -51 4628 -48 5116
rect -31 4628 -28 5116
rect -51 4622 -28 4628
rect 28 5116 51 5122
rect 28 4628 31 5116
rect 48 4628 51 5116
rect 28 4622 51 4628
rect -23 4603 23 4606
rect -23 4586 -17 4603
rect 17 4586 23 4603
rect -23 4583 23 4586
rect -23 4549 23 4552
rect -23 4532 -17 4549
rect 17 4532 23 4549
rect -23 4529 23 4532
rect -51 4507 -28 4513
rect -51 4019 -48 4507
rect -31 4019 -28 4507
rect -51 4013 -28 4019
rect 28 4507 51 4513
rect 28 4019 31 4507
rect 48 4019 51 4507
rect 28 4013 51 4019
rect -23 3994 23 3997
rect -23 3977 -17 3994
rect 17 3977 23 3994
rect -23 3974 23 3977
rect -23 3940 23 3943
rect -23 3923 -17 3940
rect 17 3923 23 3940
rect -23 3920 23 3923
rect -51 3898 -28 3904
rect -51 3410 -48 3898
rect -31 3410 -28 3898
rect -51 3404 -28 3410
rect 28 3898 51 3904
rect 28 3410 31 3898
rect 48 3410 51 3898
rect 28 3404 51 3410
rect -23 3385 23 3388
rect -23 3368 -17 3385
rect 17 3368 23 3385
rect -23 3365 23 3368
rect -23 3331 23 3334
rect -23 3314 -17 3331
rect 17 3314 23 3331
rect -23 3311 23 3314
rect -51 3289 -28 3295
rect -51 2801 -48 3289
rect -31 2801 -28 3289
rect -51 2795 -28 2801
rect 28 3289 51 3295
rect 28 2801 31 3289
rect 48 2801 51 3289
rect 28 2795 51 2801
rect -23 2776 23 2779
rect -23 2759 -17 2776
rect 17 2759 23 2776
rect -23 2756 23 2759
rect -23 2722 23 2725
rect -23 2705 -17 2722
rect 17 2705 23 2722
rect -23 2702 23 2705
rect -51 2680 -28 2686
rect -51 2192 -48 2680
rect -31 2192 -28 2680
rect -51 2186 -28 2192
rect 28 2680 51 2686
rect 28 2192 31 2680
rect 48 2192 51 2680
rect 28 2186 51 2192
rect -23 2167 23 2170
rect -23 2150 -17 2167
rect 17 2150 23 2167
rect -23 2147 23 2150
rect -23 2113 23 2116
rect -23 2096 -17 2113
rect 17 2096 23 2113
rect -23 2093 23 2096
rect -51 2071 -28 2077
rect -51 1583 -48 2071
rect -31 1583 -28 2071
rect -51 1577 -28 1583
rect 28 2071 51 2077
rect 28 1583 31 2071
rect 48 1583 51 2071
rect 28 1577 51 1583
rect -23 1558 23 1561
rect -23 1541 -17 1558
rect 17 1541 23 1558
rect -23 1538 23 1541
rect -23 1504 23 1507
rect -23 1487 -17 1504
rect 17 1487 23 1504
rect -23 1484 23 1487
rect -51 1462 -28 1468
rect -51 974 -48 1462
rect -31 974 -28 1462
rect -51 968 -28 974
rect 28 1462 51 1468
rect 28 974 31 1462
rect 48 974 51 1462
rect 28 968 51 974
rect -23 949 23 952
rect -23 932 -17 949
rect 17 932 23 949
rect -23 929 23 932
rect -23 895 23 898
rect -23 878 -17 895
rect 17 878 23 895
rect -23 875 23 878
rect -51 853 -28 859
rect -51 365 -48 853
rect -31 365 -28 853
rect -51 359 -28 365
rect 28 853 51 859
rect 28 365 31 853
rect 48 365 51 853
rect 28 359 51 365
rect -23 340 23 343
rect -23 323 -17 340
rect 17 323 23 340
rect -23 320 23 323
rect -23 286 23 289
rect -23 269 -17 286
rect 17 269 23 286
rect -23 266 23 269
rect -51 244 -28 250
rect -51 -244 -48 244
rect -31 -244 -28 244
rect -51 -250 -28 -244
rect 28 244 51 250
rect 28 -244 31 244
rect 48 -244 51 244
rect 28 -250 51 -244
rect -23 -269 23 -266
rect -23 -286 -17 -269
rect 17 -286 23 -269
rect -23 -289 23 -286
rect -23 -323 23 -320
rect -23 -340 -17 -323
rect 17 -340 23 -323
rect -23 -343 23 -340
rect -51 -365 -28 -359
rect -51 -853 -48 -365
rect -31 -853 -28 -365
rect -51 -859 -28 -853
rect 28 -365 51 -359
rect 28 -853 31 -365
rect 48 -853 51 -365
rect 28 -859 51 -853
rect -23 -878 23 -875
rect -23 -895 -17 -878
rect 17 -895 23 -878
rect -23 -898 23 -895
rect -23 -932 23 -929
rect -23 -949 -17 -932
rect 17 -949 23 -932
rect -23 -952 23 -949
rect -51 -974 -28 -968
rect -51 -1462 -48 -974
rect -31 -1462 -28 -974
rect -51 -1468 -28 -1462
rect 28 -974 51 -968
rect 28 -1462 31 -974
rect 48 -1462 51 -974
rect 28 -1468 51 -1462
rect -23 -1487 23 -1484
rect -23 -1504 -17 -1487
rect 17 -1504 23 -1487
rect -23 -1507 23 -1504
rect -23 -1541 23 -1538
rect -23 -1558 -17 -1541
rect 17 -1558 23 -1541
rect -23 -1561 23 -1558
rect -51 -1583 -28 -1577
rect -51 -2071 -48 -1583
rect -31 -2071 -28 -1583
rect -51 -2077 -28 -2071
rect 28 -1583 51 -1577
rect 28 -2071 31 -1583
rect 48 -2071 51 -1583
rect 28 -2077 51 -2071
rect -23 -2096 23 -2093
rect -23 -2113 -17 -2096
rect 17 -2113 23 -2096
rect -23 -2116 23 -2113
rect -23 -2150 23 -2147
rect -23 -2167 -17 -2150
rect 17 -2167 23 -2150
rect -23 -2170 23 -2167
rect -51 -2192 -28 -2186
rect -51 -2680 -48 -2192
rect -31 -2680 -28 -2192
rect -51 -2686 -28 -2680
rect 28 -2192 51 -2186
rect 28 -2680 31 -2192
rect 48 -2680 51 -2192
rect 28 -2686 51 -2680
rect -23 -2705 23 -2702
rect -23 -2722 -17 -2705
rect 17 -2722 23 -2705
rect -23 -2725 23 -2722
rect -23 -2759 23 -2756
rect -23 -2776 -17 -2759
rect 17 -2776 23 -2759
rect -23 -2779 23 -2776
rect -51 -2801 -28 -2795
rect -51 -3289 -48 -2801
rect -31 -3289 -28 -2801
rect -51 -3295 -28 -3289
rect 28 -2801 51 -2795
rect 28 -3289 31 -2801
rect 48 -3289 51 -2801
rect 28 -3295 51 -3289
rect -23 -3314 23 -3311
rect -23 -3331 -17 -3314
rect 17 -3331 23 -3314
rect -23 -3334 23 -3331
rect -23 -3368 23 -3365
rect -23 -3385 -17 -3368
rect 17 -3385 23 -3368
rect -23 -3388 23 -3385
rect -51 -3410 -28 -3404
rect -51 -3898 -48 -3410
rect -31 -3898 -28 -3410
rect -51 -3904 -28 -3898
rect 28 -3410 51 -3404
rect 28 -3898 31 -3410
rect 48 -3898 51 -3410
rect 28 -3904 51 -3898
rect -23 -3923 23 -3920
rect -23 -3940 -17 -3923
rect 17 -3940 23 -3923
rect -23 -3943 23 -3940
rect -23 -3977 23 -3974
rect -23 -3994 -17 -3977
rect 17 -3994 23 -3977
rect -23 -3997 23 -3994
rect -51 -4019 -28 -4013
rect -51 -4507 -48 -4019
rect -31 -4507 -28 -4019
rect -51 -4513 -28 -4507
rect 28 -4019 51 -4013
rect 28 -4507 31 -4019
rect 48 -4507 51 -4019
rect 28 -4513 51 -4507
rect -23 -4532 23 -4529
rect -23 -4549 -17 -4532
rect 17 -4549 23 -4532
rect -23 -4552 23 -4549
rect -23 -4586 23 -4583
rect -23 -4603 -17 -4586
rect 17 -4603 23 -4586
rect -23 -4606 23 -4603
rect -51 -4628 -28 -4622
rect -51 -5116 -48 -4628
rect -31 -5116 -28 -4628
rect -51 -5122 -28 -5116
rect 28 -4628 51 -4622
rect 28 -5116 31 -4628
rect 48 -5116 51 -4628
rect 28 -5122 51 -5116
rect -23 -5141 23 -5138
rect -23 -5158 -17 -5141
rect 17 -5158 23 -5141
rect -23 -5161 23 -5158
rect -23 -5195 23 -5192
rect -23 -5212 -17 -5195
rect 17 -5212 23 -5195
rect -23 -5215 23 -5212
rect -51 -5237 -28 -5231
rect -51 -5725 -48 -5237
rect -31 -5725 -28 -5237
rect -51 -5731 -28 -5725
rect 28 -5237 51 -5231
rect 28 -5725 31 -5237
rect 48 -5725 51 -5237
rect 28 -5731 51 -5725
rect -23 -5750 23 -5747
rect -23 -5767 -17 -5750
rect 17 -5767 23 -5750
rect -23 -5770 23 -5767
<< properties >>
string FIXED_BBOX -96 -5809 96 5809
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.5 m 19 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
