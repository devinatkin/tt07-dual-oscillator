** sch_path: /home/dmatkin/tt07-dual-oscillator/xschem/oscillator_21MHZ.sch
.subckt oscillator_21MHZ VCC OUT VSS
*.PININFO VCC:B VSS:B OUT:O
x1[20] INI[19] OUT_INI VCC VSS inverter
x1[19] INI[18] INI[19] VCC VSS inverter
x1[18] INI[17] INI[18] VCC VSS inverter
x1[17] INI[16] INI[17] VCC VSS inverter
x1[16] INI[15] INI[16] VCC VSS inverter
x1[15] INI[14] INI[15] VCC VSS inverter
x1[14] INI[13] INI[14] VCC VSS inverter
x1[13] INI[12] INI[13] VCC VSS inverter
x1[12] INI[11] INI[12] VCC VSS inverter
x1[11] INI[10] INI[11] VCC VSS inverter
x1[10] INI[9] INI[10] VCC VSS inverter
x1[9] INI[8] INI[9] VCC VSS inverter
x1[8] INI[7] INI[8] VCC VSS inverter
x1[7] INI[6] INI[7] VCC VSS inverter
x1[6] INI[5] INI[6] VCC VSS inverter
x1[5] INI[4] INI[5] VCC VSS inverter
x1[4] INI[3] INI[4] VCC VSS inverter
x1[3] INI[2] INI[3] VCC VSS inverter
x1[2] INI[1] INI[2] VCC VSS inverter
x1[1] INI[0] INI[1] VCC VSS inverter
x1[0] OUT_INI INI[0] VCC VSS inverter
x1 OUT OUT_INI VCC VSS inverter
.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/dmatkin/tt07-dual-oscillator/xschem/inverter.sym
** sch_path: /home/dmatkin/tt07-dual-oscillator/xschem/inverter.sch
.subckt inverter OUT IN VCC VSS
*.PININFO VCC:B VSS:B IN:I OUT:O
XM1 OUT IN net1 VCC sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 m=1
XM2 OUT IN net2 VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM3 net1 VSS VCC VCC sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 m=1
XM4 net2 VCC VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
.ends

.end
