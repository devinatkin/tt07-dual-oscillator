magic
tech sky130A
magscale 1 2
timestamp 1715270440
<< metal1 >>
rect 7156 28339 7284 28673
rect 7614 28339 7620 28673
rect 6331 8875 6531 10333
rect 4577 1194 4782 2655
rect 6332 1857 6530 8875
rect 6332 1659 27768 1857
rect 26871 1325 27041 1659
rect 4577 989 26379 1194
rect 26865 1155 26871 1325
rect 27041 1155 27047 1325
rect 31264 1193 31469 1199
rect 26174 804 26379 989
rect 27468 988 31264 1193
rect 27468 804 27673 988
rect 31264 982 31469 988
rect 26174 599 27673 804
<< via1 >>
rect 5406 28462 5720 28662
rect 7284 28339 7614 28673
rect 26871 1155 27041 1325
rect 31264 988 31469 1193
<< metal2 >>
rect 1214 29124 1223 29483
rect 1582 29124 5745 29483
rect 5386 28662 5745 29124
rect 5386 28462 5406 28662
rect 5720 28462 5745 28662
rect 5386 28446 5745 28462
rect 7284 28673 7614 28679
rect 7614 28341 8029 28671
rect 8359 28341 8368 28671
rect 7284 28333 7614 28339
rect 26871 1325 27041 1331
rect 31264 1193 31469 1202
rect 26871 1126 27041 1155
rect 26867 966 26876 1126
rect 27036 966 27045 1126
rect 31258 988 31264 1193
rect 31469 988 31475 1193
rect 31264 979 31469 988
rect 26871 961 27041 966
<< via2 >>
rect 1223 29124 1582 29483
rect 8029 28341 8359 28671
rect 26876 966 27036 1126
rect 31264 988 31469 1193
<< metal3 >>
rect 1212 29119 1218 29488
rect 1577 29483 1587 29488
rect 1582 29124 1587 29483
rect 1577 29119 1587 29124
rect 8024 28671 8364 28676
rect 8024 28341 8029 28671
rect 8359 28341 8805 28671
rect 9135 28341 9141 28671
rect 8024 28336 8364 28341
rect 31259 1193 31474 1198
rect 26871 1126 27041 1131
rect 26871 966 26876 1126
rect 27036 966 27041 1126
rect 31259 988 31264 1193
rect 31469 988 31474 1193
rect 31259 983 31474 988
rect 26871 522 27041 966
rect 31264 881 31469 983
rect 31264 670 31469 676
rect 26866 354 26872 522
rect 27040 354 27046 522
rect 26871 353 27041 354
rect 31293 65 31440 670
<< via3 >>
rect 1218 29483 1577 29488
rect 1218 29124 1223 29483
rect 1223 29124 1577 29483
rect 1218 29119 1577 29124
rect 8805 28341 9135 28671
rect 31264 676 31469 881
rect 26872 354 27040 522
<< metal4 >>
rect 798 44644 858 45152
rect 1534 44644 1594 45152
rect 2270 44644 2330 45152
rect 3006 44644 3066 45152
rect 3742 44644 3802 45152
rect 4478 44644 4538 45152
rect 5214 44644 5274 45152
rect 5950 44644 6010 45152
rect 6686 44644 6746 45152
rect 7422 44644 7482 45152
rect 8158 44644 8218 45152
rect 8894 44644 8954 45152
rect 9630 44644 9690 45152
rect 10366 44644 10426 45152
rect 11102 44644 11162 45152
rect 11838 44644 11898 45152
rect 12574 44644 12634 45152
rect 13310 44644 13370 45152
rect 14046 44644 14106 45152
rect 14782 44644 14842 45152
rect 15518 44644 15578 45152
rect 16254 44644 16314 45152
rect 16990 44644 17050 45152
rect 17726 44644 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 594 44324 17918 44644
rect 200 29483 500 44152
rect 1217 29488 1578 29489
rect 1217 29483 1218 29488
rect 200 29124 1218 29483
rect 200 1000 500 29124
rect 1217 29119 1218 29124
rect 1577 29119 1578 29488
rect 1217 29118 1578 29119
rect 8804 28671 9136 28672
rect 9800 28671 10100 44324
rect 8804 28341 8805 28671
rect 9135 28341 10100 28671
rect 8804 28340 9136 28341
rect 9800 1000 10100 28341
rect 31263 881 31470 882
rect 31263 676 31264 881
rect 31469 676 31470 881
rect 31263 675 31470 676
rect 26871 522 27041 523
rect 26871 354 26872 522
rect 27040 354 27041 522
rect 26871 200 27041 354
rect 31307 200 31426 675
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 200
use top  top_0 ~/tt07-dual-oscillator/mag
timestamp 1715268526
transform 0 1 7644 -1 0 29078
box 404 -3722 26563 -430
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
