magic
tech sky130A
timestamp 1716524512
<< pwell >>
rect -191 -152 1172 1465
<< psubdiff >>
rect -156 1417 -121 1434
rect 1099 1417 1130 1434
rect -156 1393 -139 1417
rect -156 -105 -139 -68
rect 1113 1384 1130 1417
rect 1113 -105 1130 -77
rect -156 -122 -94 -105
rect 1034 -122 1130 -105
<< psubdiffcont >>
rect -121 1417 1099 1434
rect -156 -68 -139 1393
rect 1113 -77 1130 1384
rect -94 -122 1034 -105
<< locali >>
rect -156 1417 -121 1434
rect 1099 1417 1130 1434
rect -156 1393 -139 1417
rect -156 -105 -139 -68
rect 1113 1384 1130 1417
rect 1113 -105 1130 -77
rect -156 -122 -94 -105
rect 1034 -122 1130 -105
<< viali >>
rect -93 -122 128 -105
<< metal1 >>
rect 29 1348 730 1349
rect 28 1346 730 1348
rect 28 1319 431 1346
rect 522 1319 730 1346
rect 28 1317 730 1319
rect 28 1269 129 1317
rect 408 1316 571 1317
rect 48 1262 129 1269
rect 629 1263 730 1317
rect -11 1069 -1 1241
rect 27 1069 31 1241
rect 134 1214 223 1246
rect 134 1099 147 1214
rect 203 1099 223 1214
rect 134 741 223 1099
rect 591 1242 653 1245
rect 591 1059 596 1242
rect 629 1059 653 1242
rect 591 1056 653 1059
rect 734 1214 823 1247
rect 734 1099 748 1214
rect 804 1099 823 1214
rect 335 1004 388 1013
rect 335 852 346 1004
rect 380 852 388 1004
rect 335 840 388 852
rect 734 742 823 1099
rect 936 1001 989 1013
rect 936 851 939 1001
rect 984 851 989 1001
rect 936 840 989 851
rect 229 650 329 724
rect 827 651 929 725
rect 574 650 929 651
rect 31 649 929 650
rect 30 618 929 649
rect 30 563 131 618
rect 574 617 929 618
rect 422 590 525 599
rect 422 588 435 590
rect 228 563 435 588
rect 519 563 525 590
rect 33 561 129 563
rect 228 560 525 563
rect 627 560 732 617
rect 825 588 929 594
rect 825 562 837 588
rect 921 562 929 588
rect 825 559 929 562
rect 135 546 205 547
rect -7 492 45 501
rect -7 359 0 492
rect 31 359 45 492
rect -7 349 45 359
rect 135 176 224 546
rect 590 492 642 502
rect 590 359 605 492
rect 636 359 642 492
rect 590 350 642 359
rect 135 61 152 176
rect 208 61 224 176
rect 323 282 375 292
rect 323 149 333 282
rect 364 149 375 282
rect 323 140 375 149
rect 734 181 823 523
rect 135 42 224 61
rect 734 66 753 181
rect 809 66 823 181
rect 922 281 974 295
rect 922 148 934 281
rect 965 148 974 281
rect 922 143 974 148
rect 734 41 823 66
rect -113 -105 138 -83
rect -113 -122 -93 -105
rect 128 -122 138 -105
rect -113 -141 138 -122
<< via1 >>
rect 431 1319 522 1346
rect -1 1069 27 1241
rect 147 1099 203 1214
rect 596 1059 629 1242
rect 748 1099 804 1214
rect 346 852 380 1004
rect 939 851 984 1001
rect 435 563 519 590
rect 837 562 921 588
rect 0 359 31 492
rect 605 359 636 492
rect 152 61 208 176
rect 333 149 364 282
rect 753 66 809 181
rect 934 148 965 281
<< metal2 >>
rect 427 1346 525 1349
rect 427 1319 431 1346
rect 522 1319 525 1346
rect 427 1286 525 1319
rect -11 1241 32 1248
rect -11 1238 -1 1241
rect 27 1238 32 1241
rect -11 1062 -6 1238
rect 29 1062 32 1238
rect -11 1056 32 1062
rect 134 1214 223 1246
rect 134 1099 147 1214
rect 203 1099 223 1214
rect 134 802 223 1099
rect 133 791 223 802
rect 133 746 138 791
rect 217 746 223 791
rect -6 492 42 497
rect -6 359 0 492
rect 31 486 42 492
rect 39 362 42 486
rect 133 404 223 746
rect 323 1005 390 1013
rect 323 847 344 1005
rect 379 1004 390 1005
rect 380 852 390 1004
rect 379 847 390 852
rect 323 658 390 847
rect 427 729 524 1286
rect 549 1245 649 1246
rect 549 1242 653 1245
rect 549 1234 596 1242
rect 542 1059 596 1234
rect 629 1059 653 1242
rect 542 1056 653 1059
rect 735 1214 825 1241
rect 735 1099 748 1214
rect 804 1099 825 1214
rect 542 1053 649 1056
rect 427 679 525 729
rect 31 359 42 362
rect -6 351 42 359
rect 134 176 223 404
rect 324 486 388 658
rect 428 592 525 679
rect 428 563 434 592
rect 519 563 525 592
rect 428 542 525 563
rect 324 360 333 486
rect 381 360 388 486
rect 324 356 388 360
rect 134 93 152 176
rect 208 93 223 176
rect 325 284 373 288
rect 542 284 579 1053
rect 735 876 825 1099
rect 732 794 825 876
rect 935 1002 990 1013
rect 935 1001 944 1002
rect 979 1001 990 1002
rect 935 851 939 1001
rect 984 851 990 1001
rect 935 844 944 851
rect 979 844 990 851
rect 935 840 990 844
rect 732 744 742 794
rect 820 744 825 794
rect 732 743 825 744
rect 732 539 798 743
rect 828 591 929 595
rect 828 559 834 591
rect 924 559 929 591
rect 828 552 929 559
rect 595 492 643 500
rect 595 490 605 492
rect 636 490 643 492
rect 595 366 601 490
rect 640 366 643 490
rect 595 359 605 366
rect 636 359 643 366
rect 595 354 643 359
rect 325 145 330 284
rect 365 145 373 284
rect 530 272 588 284
rect 530 159 534 272
rect 584 159 588 272
rect 530 149 588 159
rect 732 181 822 539
rect 325 142 373 145
rect 134 46 143 93
rect 215 46 223 93
rect 134 42 223 46
rect 732 95 753 181
rect 809 95 822 181
rect 926 282 974 290
rect 926 148 934 282
rect 964 281 974 282
rect 965 148 974 281
rect 926 144 974 148
rect 732 48 745 95
rect 817 48 822 95
rect 732 41 822 48
<< via2 >>
rect -6 1069 -1 1238
rect -1 1069 27 1238
rect 27 1069 29 1238
rect -6 1062 29 1069
rect 138 746 217 791
rect 0 362 31 486
rect 31 362 39 486
rect 344 1004 379 1005
rect 344 852 346 1004
rect 346 852 379 1004
rect 344 847 379 852
rect 598 1060 628 1237
rect 434 590 519 592
rect 434 563 435 590
rect 435 563 519 590
rect 333 360 381 486
rect 944 1001 979 1002
rect 944 851 979 1001
rect 944 844 979 851
rect 742 744 820 794
rect 834 588 924 591
rect 834 562 837 588
rect 837 562 921 588
rect 921 562 924 588
rect 834 559 924 562
rect 601 366 605 490
rect 605 366 636 490
rect 636 366 640 490
rect 330 282 365 284
rect 330 149 333 282
rect 333 149 364 282
rect 364 149 365 282
rect 330 145 365 149
rect 534 159 584 272
rect 143 61 152 93
rect 152 61 208 93
rect 208 61 215 93
rect 143 46 215 61
rect 934 281 964 282
rect 934 149 964 281
rect 745 66 753 95
rect 753 66 809 95
rect 809 66 817 95
rect 745 48 817 66
<< metal3 >>
rect -22 1238 632 1247
rect -22 1062 -6 1238
rect 29 1237 632 1238
rect 29 1062 598 1237
rect -22 1060 598 1062
rect 628 1060 632 1237
rect -22 1056 632 1060
rect -22 1055 86 1056
rect 335 1005 991 1014
rect 335 847 344 1005
rect 379 1002 991 1005
rect 379 847 944 1002
rect 335 844 944 847
rect 979 844 991 1002
rect 335 839 991 844
rect 134 794 823 797
rect 134 791 742 794
rect 134 746 138 791
rect 217 746 742 791
rect 134 744 742 746
rect 820 744 823 794
rect 134 740 823 744
rect 428 592 929 595
rect 428 563 434 592
rect 519 591 929 592
rect 519 563 834 591
rect 428 559 834 563
rect 924 559 929 591
rect 428 542 929 559
rect -8 494 101 495
rect -8 490 667 494
rect -8 486 601 490
rect -8 362 0 486
rect 39 362 333 486
rect -8 360 333 362
rect 381 366 601 486
rect 640 366 667 490
rect 381 360 667 366
rect -8 358 667 360
rect -8 357 626 358
rect -8 356 101 357
rect 316 285 378 295
rect 316 284 447 285
rect 316 145 330 284
rect 365 283 447 284
rect 916 283 978 294
rect 365 282 1004 283
rect 365 272 934 282
rect 365 159 534 272
rect 584 159 934 272
rect 365 149 934 159
rect 964 149 1004 282
rect 365 146 1004 149
rect 365 145 447 146
rect 894 145 1004 146
rect 316 134 378 145
rect 916 135 978 145
rect 133 95 822 99
rect 133 93 745 95
rect 133 46 143 93
rect 215 48 745 93
rect 817 48 822 95
rect 215 46 822 48
rect 133 42 822 46
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_0
timestamp 1716523272
transform 1 0 879 0 1 994
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_1
timestamp 1716523272
transform 1 0 79 0 1 294
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_2
timestamp 1716523272
transform 1 0 279 0 1 294
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_3
timestamp 1716523272
transform 1 0 679 0 1 294
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_4
timestamp 1716523272
transform 1 0 879 0 1 294
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_5
timestamp 1716523272
transform 1 0 79 0 1 994
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_6
timestamp 1716523272
transform 1 0 279 0 1 994
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_7
timestamp 1716523272
transform 1 0 679 0 1 994
box -79 -294 79 294
<< labels >>
flabel metal1 -113 -105 138 -83 0 FreeSans 240 0 0 0 VSS
port 1 nsew
flabel metal3 215 42 745 99 0 FreeSans 240 0 0 0 S
port 2 nsew
flabel metal1 29 1317 431 1349 0 FreeSans 240 0 0 0 INA
port 3 nsew
flabel metal1 574 617 929 651 0 FreeSans 240 0 0 0 INB
port 4 nsew
flabel metal3 29 1056 598 1247 0 FreeSans 240 0 0 0 DA
port 5 nsew
flabel metal3 381 357 601 494 0 FreeSans 240 0 0 0 DB
port 6 nsew
<< end >>
