magic
tech sky130A
magscale 1 2
timestamp 1716849570
<< nwell >>
rect -246 -969 246 969
<< pmoslvt >>
rect -50 -750 50 750
<< pdiff >>
rect -108 738 -50 750
rect -108 -738 -96 738
rect -62 -738 -50 738
rect -108 -750 -50 -738
rect 50 738 108 750
rect 50 -738 62 738
rect 96 -738 108 738
rect 50 -750 108 -738
<< pdiffc >>
rect -96 -738 -62 738
rect 62 -738 96 738
<< nsubdiff >>
rect -210 899 -114 933
rect 114 899 210 933
rect -210 837 -176 899
rect 176 837 210 899
rect -210 -899 -176 -837
rect 176 -899 210 -837
rect -210 -933 -114 -899
rect 114 -933 210 -899
<< nsubdiffcont >>
rect -114 899 114 933
rect -210 -837 -176 837
rect 176 -837 210 837
rect -114 -933 114 -899
<< poly >>
rect -50 831 50 847
rect -50 797 -34 831
rect 34 797 50 831
rect -50 750 50 797
rect -50 -797 50 -750
rect -50 -831 -34 -797
rect 34 -831 50 -797
rect -50 -847 50 -831
<< polycont >>
rect -34 797 34 831
rect -34 -831 34 -797
<< locali >>
rect -210 899 -114 933
rect 114 899 210 933
rect -210 837 -176 899
rect 176 837 210 899
rect -50 797 -34 831
rect 34 797 50 831
rect -96 738 -62 754
rect -96 -754 -62 -738
rect 62 738 96 754
rect 62 -754 96 -738
rect -50 -831 -34 -797
rect 34 -831 50 -797
rect -210 -899 -176 -837
rect 176 -899 210 -837
rect -210 -933 -114 -899
rect 114 -933 210 -899
<< viali >>
rect -34 797 34 831
rect -96 -738 -62 738
rect 62 -738 96 738
rect -34 -831 34 -797
<< metal1 >>
rect -46 831 46 837
rect -46 797 -34 831
rect 34 797 46 831
rect -46 791 46 797
rect -102 738 -56 750
rect -102 -738 -96 738
rect -62 -738 -56 738
rect -102 -750 -56 -738
rect 56 738 102 750
rect 56 -738 62 738
rect 96 -738 102 738
rect 56 -750 102 -738
rect -46 -797 46 -791
rect -46 -831 -34 -797
rect 34 -831 46 -797
rect -46 -837 46 -831
<< properties >>
string FIXED_BBOX -193 -916 193 916
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 7.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
