magic
tech sky130A
timestamp 1717178954
<< nwell >>
rect 2611 240 4338 630
rect 4325 239 4338 240
<< pwell >>
rect 1933 1225 4337 2936
rect 1934 631 4337 1225
rect 2180 630 4337 631
<< metal1 >>
rect 1749 2847 2033 2904
rect 1934 2057 2033 2847
rect 1898 2001 2033 2057
rect 919 1962 2033 2001
rect 1898 1934 2033 1962
rect 1631 1563 1713 1578
rect 1631 1421 1644 1563
rect 1702 1421 1713 1563
rect 1631 1398 1713 1421
rect 1010 1306 1017 1354
rect 1094 1306 1099 1354
rect 1010 1294 1099 1306
rect 790 1173 925 1188
rect 790 1095 809 1173
rect 900 1095 925 1173
rect 790 1077 925 1095
rect 1934 611 2033 1934
rect 2604 540 2740 630
rect 1600 473 1733 488
rect 1600 388 1616 473
rect 1713 388 1733 473
rect 1600 377 1733 388
rect 2657 180 2740 540
rect 649 -1261 735 -323
rect 2712 -417 2862 -399
rect 2712 -509 2723 -417
rect 2846 -509 2862 -417
rect 2712 -517 2862 -509
rect 2394 -598 2840 -586
rect 2394 -659 2412 -598
rect 2494 -659 2840 -598
rect 2394 -673 2840 -659
rect 1724 -1061 1821 -1057
rect 819 -1099 1821 -1061
rect 819 -1100 1734 -1099
rect 1724 -1162 1734 -1100
rect 1815 -1162 1821 -1099
rect 1724 -1172 1821 -1162
rect 1887 -1259 1988 -1253
rect 1767 -1296 1988 -1259
rect 1767 -1302 1965 -1296
rect 2571 -1302 2722 -1266
<< via1 >>
rect 1644 1421 1702 1563
rect 1017 1306 1094 1355
rect 809 1095 900 1173
rect 1616 388 1713 473
rect 2723 -509 2846 -417
rect 2412 -659 2494 -598
rect 1734 -1162 1815 -1099
rect 2063 -1240 2089 -1111
<< metal2 >>
rect 1643 1579 1716 1886
rect 1585 1563 1716 1579
rect 1585 1421 1644 1563
rect 1702 1421 1716 1563
rect 1010 1355 1099 1360
rect 1010 1306 1017 1355
rect 1094 1306 1099 1355
rect 790 1173 925 1188
rect 790 1095 809 1173
rect 900 1095 925 1173
rect 790 1077 925 1095
rect 1010 989 1099 1306
rect 1585 1147 1716 1421
rect 1890 1304 2083 1305
rect 1890 1284 2124 1304
rect 1585 1083 1855 1147
rect 1585 1082 1716 1083
rect 1010 836 1021 989
rect 1085 836 1099 989
rect 1010 821 1099 836
rect 1798 720 1855 1083
rect 1890 879 1913 1284
rect 2080 879 2124 1284
rect 1890 858 2124 879
rect 1890 850 2182 858
rect 1798 606 1807 720
rect 1842 606 1855 720
rect 1600 475 1733 488
rect 1600 473 1650 475
rect 1600 388 1616 473
rect 1720 410 1733 475
rect 1713 388 1733 410
rect 1600 377 1733 388
rect 1798 264 1855 606
rect 2053 690 2182 850
rect 1798 243 1889 264
rect 1798 136 1814 243
rect 1865 136 1889 243
rect 1798 118 1889 136
rect 1381 -147 1468 -141
rect 1381 -192 1392 -147
rect 1462 -192 1468 -147
rect 1381 -548 1468 -192
rect 1799 -436 1889 118
rect 2053 -256 2124 690
rect 2341 678 2597 689
rect 2341 632 2371 678
rect 2553 632 2597 678
rect 2341 378 2597 632
rect 2331 267 2468 278
rect 2331 164 2349 267
rect 2453 164 2468 267
rect 2331 -214 2468 164
rect 2053 -355 2067 -256
rect 2112 -355 2124 -256
rect 2053 -376 2124 -355
rect 1799 -497 1809 -436
rect 1879 -497 1889 -436
rect 1799 -504 1889 -497
rect 2712 -417 2862 -399
rect 2712 -509 2723 -417
rect 2846 -509 2862 -417
rect 2712 -517 2862 -509
rect 1381 -629 1389 -548
rect 1455 -629 1468 -548
rect 1381 -634 1468 -629
rect 2393 -598 2517 -586
rect 2393 -659 2412 -598
rect 2494 -659 2517 -598
rect 1723 -1099 1870 -1060
rect 1723 -1201 1734 -1099
rect 1815 -1101 1870 -1099
rect 1854 -1201 1870 -1101
rect 1723 -1207 1870 -1201
rect 2031 -1101 2135 -1095
rect 2031 -1198 2038 -1101
rect 2126 -1198 2135 -1101
rect 2031 -1240 2063 -1198
rect 2089 -1240 2135 -1198
rect 2393 -1100 2517 -659
rect 2393 -1196 2408 -1100
rect 2500 -1196 2517 -1100
rect 2393 -1209 2517 -1196
rect 2031 -1253 2135 -1240
<< via2 >>
rect 809 1095 900 1173
rect 1021 836 1085 989
rect 1913 879 2080 1284
rect 1807 606 1842 720
rect 1650 473 1720 475
rect 1650 410 1713 473
rect 1713 410 1720 473
rect 1814 136 1865 243
rect 1392 -192 1462 -147
rect 2371 632 2553 678
rect 2349 164 2453 267
rect 2067 -355 2112 -256
rect 1809 -497 1879 -436
rect 2723 -509 2846 -417
rect 1389 -629 1455 -548
rect 1734 -1162 1815 -1101
rect 1815 -1162 1854 -1101
rect 1734 -1201 1854 -1162
rect 2038 -1111 2126 -1101
rect 2038 -1198 2063 -1111
rect 2063 -1198 2089 -1111
rect 2089 -1198 2126 -1111
rect 2408 -1196 2500 -1100
<< metal3 >>
rect 1890 1286 2143 1309
rect 790 1173 925 1188
rect 790 1095 809 1173
rect 900 1095 925 1173
rect 790 1077 925 1095
rect 1890 875 1904 1286
rect 2082 936 2143 1286
rect 2082 875 2138 936
rect 1890 850 2138 875
rect 1783 720 2015 727
rect 1783 606 1807 720
rect 1842 692 2015 720
rect 1842 691 2038 692
rect 1842 689 2195 691
rect 1842 678 2597 689
rect 1842 632 2371 678
rect 2553 632 2597 678
rect 1842 606 2597 632
rect 1783 600 2597 606
rect 1633 475 1766 509
rect 1633 410 1650 475
rect 1720 410 1766 475
rect 1633 398 1766 410
rect 2332 294 2896 310
rect 2332 267 2788 294
rect 1211 243 1878 254
rect 1211 136 1814 243
rect 1865 136 1878 243
rect 2332 164 2349 267
rect 2453 179 2788 267
rect 2876 179 2896 294
rect 2453 164 2896 179
rect 2332 156 2896 164
rect 1211 117 1878 136
rect 2048 -256 2849 -239
rect 2048 -355 2067 -256
rect 2112 -355 2849 -256
rect 2048 -375 2849 -355
rect 3879 -367 3981 -241
rect 2707 -417 2857 -409
rect 2707 -425 2723 -417
rect 1799 -436 2723 -425
rect 1799 -497 1809 -436
rect 1879 -497 2723 -436
rect 1799 -504 2723 -497
rect 2707 -509 2723 -504
rect 2846 -509 2857 -417
rect 2707 -527 2857 -509
rect 1723 -1100 2516 -1092
rect 1723 -1101 2408 -1100
rect 1723 -1201 1734 -1101
rect 1854 -1198 2038 -1101
rect 2126 -1196 2408 -1101
rect 2500 -1196 2516 -1100
rect 2126 -1198 2516 -1196
rect 1854 -1201 2516 -1198
rect 1723 -1208 2516 -1201
<< via3 >>
rect 1904 1284 2082 1286
rect 1904 879 1913 1284
rect 1913 879 2080 1284
rect 2080 879 2082 1284
rect 1904 875 2082 879
rect 2788 179 2876 294
<< metal4 >>
rect 2086 1305 2152 2157
rect 1885 1286 2152 1305
rect 1885 875 1904 1286
rect 2082 936 2152 1286
rect 2082 875 2138 936
rect 1885 850 2138 875
rect 2270 859 4232 2121
rect 2768 567 3047 859
rect 2770 294 2892 567
rect 2770 179 2788 294
rect 2876 179 2892 294
rect 2770 161 2892 179
use active-resistor  active-resistor_0
timestamp 1717178954
transform 1 0 209 0 1 -422
box 1725 -892 2402 1053
use activeload  activeload_0
timestamp 1717178954
transform 1 0 546 0 1 1226
box 0 0 1387 1710
use indiff  indiff_0
timestamp 1717178954
transform 1 0 762 0 1 -240
box -191 -152 1172 1465
use second_stage  second_stage_0
timestamp 1717178954
transform 1 0 2725 0 1 -1233
box -114 -82 1613 1473
use sky130_fd_pr__cap_mim_m3_1_NY928X  sky130_fd_pr__cap_mim_m3_1_NY928X_0
timestamp 1717178954
transform -1 0 3178 0 -1 1490
box -1093 -670 1093 670
use tail_current  tail_current_0
timestamp 1717178954
transform 1 0 546 0 1 -1314
box 0 0 1387 922
<< labels >>
flabel metal1 819 -1100 1821 -1061 0 FreeSans 400 0 0 0 IBIAS
port 0 nsew
flabel metal3 1720 398 1766 509 0 FreeSans 400 0 0 0 INB
port 1 nsew
flabel metal3 900 1077 925 1188 0 FreeSans 400 0 0 0 INA
port 2 nsew
flabel space 1754 -1296 2000 -1253 0 FreeSans 320 0 0 0 VSS
port 3 nsew
flabel metal1 1910 2847 2019 2904 0 FreeSans 320 0 0 0 VCC
port 4 nsew
flabel metal3 3879 -367 3981 -241 0 FreeSans 320 0 0 0 OUT
port 5 nsew
flabel metal1 1767 -1302 1965 -1259 0 FreeSans 160 0 0 0 VSS
port 6 nsew
<< end >>
