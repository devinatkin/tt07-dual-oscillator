magic
tech sky130A
magscale 1 2
timestamp 1716506474
<< pwell >>
rect -739 -1082 739 1082
<< psubdiff >>
rect -703 1012 -607 1046
rect 607 1012 703 1046
rect -703 950 -669 1012
rect 669 950 703 1012
rect -703 -1012 -669 -950
rect 669 -1012 703 -950
rect -703 -1046 -607 -1012
rect 607 -1046 703 -1012
<< psubdiffcont >>
rect -607 1012 607 1046
rect -703 -950 -669 950
rect 669 -950 703 950
rect -607 -1046 607 -1012
<< xpolycontact >>
rect -573 484 573 916
rect -573 -916 573 -484
<< xpolyres >>
rect -573 -484 573 484
<< locali >>
rect -703 1012 -607 1046
rect 607 1012 703 1046
rect -703 950 -669 1012
rect 669 950 703 1012
rect -703 -1012 -669 -950
rect 669 -1012 703 -950
rect -703 -1046 -607 -1012
rect 607 -1046 703 -1012
<< viali >>
rect -557 501 557 898
rect -557 -898 557 -501
<< metal1 >>
rect -569 898 569 904
rect -569 501 -557 898
rect 557 501 569 898
rect -569 495 569 501
rect -569 -501 569 -495
rect -569 -898 -557 -501
rect 557 -898 569 -501
rect -569 -904 569 -898
<< properties >>
string FIXED_BBOX -686 -1029 686 1029
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 5.730 l 5 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 1.81k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
