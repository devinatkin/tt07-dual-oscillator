VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_devinatkin_dual_oscillator
  CLASS BLOCK ;
  FOREIGN tt_um_devinatkin_dual_oscillator ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 533.479614 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 14.250 9.990 17.450 221.590 ;
      LAYER pwell ;
        RECT 17.450 220.890 20.740 221.590 ;
        RECT 20.960 220.950 24.250 221.650 ;
        RECT 17.450 10.620 20.750 220.890 ;
        RECT 20.950 10.620 24.250 220.950 ;
        RECT 17.450 9.970 20.740 10.620 ;
        RECT 20.960 9.970 24.250 10.620 ;
      LAYER nwell ;
        RECT 24.250 9.990 27.450 221.650 ;
      LAYER li1 ;
        RECT 14.430 220.490 17.260 220.540 ;
        RECT 14.310 220.370 17.260 220.490 ;
        RECT 14.310 218.960 14.600 220.370 ;
        RECT 14.940 219.500 15.110 219.830 ;
        RECT 15.325 219.800 16.365 219.970 ;
        RECT 15.325 219.360 16.365 219.530 ;
        RECT 16.580 219.500 16.750 219.830 ;
        RECT 17.090 218.960 17.260 220.370 ;
        RECT 14.310 218.840 17.260 218.960 ;
        RECT 14.430 218.790 17.260 218.840 ;
        RECT 17.820 220.460 20.560 220.530 ;
        RECT 21.140 220.520 23.880 220.590 ;
        RECT 17.820 220.360 20.690 220.460 ;
        RECT 17.820 218.950 17.990 220.360 ;
        RECT 18.330 219.490 18.500 219.820 ;
        RECT 18.670 219.790 19.710 219.960 ;
        RECT 18.670 219.350 19.710 219.520 ;
        RECT 19.880 219.490 20.050 219.820 ;
        RECT 20.390 218.950 20.690 220.360 ;
        RECT 17.820 218.810 20.690 218.950 ;
        RECT 21.010 220.420 23.880 220.520 ;
        RECT 21.010 219.010 21.310 220.420 ;
        RECT 21.650 219.550 21.820 219.880 ;
        RECT 21.990 219.850 23.030 220.020 ;
        RECT 21.990 219.410 23.030 219.580 ;
        RECT 23.200 219.550 23.370 219.880 ;
        RECT 23.710 219.010 23.880 220.420 ;
        RECT 21.010 218.870 23.880 219.010 ;
        RECT 24.440 220.550 27.270 220.600 ;
        RECT 24.440 220.430 27.390 220.550 ;
        RECT 24.440 219.020 24.610 220.430 ;
        RECT 24.950 219.560 25.120 219.890 ;
        RECT 25.335 219.860 26.375 220.030 ;
        RECT 25.335 219.420 26.375 219.590 ;
        RECT 26.590 219.560 26.760 219.890 ;
        RECT 27.100 219.020 27.390 220.430 ;
        RECT 24.440 218.940 27.390 219.020 ;
        RECT 17.820 218.780 20.560 218.810 ;
        RECT 14.430 218.390 17.260 218.440 ;
        RECT 14.310 218.270 17.260 218.390 ;
        RECT 14.310 216.860 14.600 218.270 ;
        RECT 14.940 217.400 15.110 217.730 ;
        RECT 15.325 217.700 16.365 217.870 ;
        RECT 15.325 217.260 16.365 217.430 ;
        RECT 16.580 217.400 16.750 217.730 ;
        RECT 17.090 216.860 17.260 218.270 ;
        RECT 14.310 216.740 17.260 216.860 ;
        RECT 14.430 216.690 17.260 216.740 ;
        RECT 17.820 218.360 20.560 218.430 ;
        RECT 21.140 218.420 23.880 218.870 ;
        RECT 17.820 218.260 20.690 218.360 ;
        RECT 17.820 216.850 17.990 218.260 ;
        RECT 18.330 217.390 18.500 217.720 ;
        RECT 18.670 217.690 19.710 217.860 ;
        RECT 18.670 217.250 19.710 217.420 ;
        RECT 19.880 217.390 20.050 217.720 ;
        RECT 20.390 216.850 20.690 218.260 ;
        RECT 17.820 216.710 20.690 216.850 ;
        RECT 21.010 218.320 23.880 218.420 ;
        RECT 24.430 218.330 27.390 218.940 ;
        RECT 21.010 216.910 21.310 218.320 ;
        RECT 21.650 217.450 21.820 217.780 ;
        RECT 21.990 217.750 23.030 217.920 ;
        RECT 21.990 217.310 23.030 217.480 ;
        RECT 23.200 217.450 23.370 217.780 ;
        RECT 23.710 216.910 23.880 218.320 ;
        RECT 21.010 216.770 23.880 216.910 ;
        RECT 24.440 216.920 24.610 218.330 ;
        RECT 24.950 217.460 25.120 217.790 ;
        RECT 25.335 217.760 26.375 217.930 ;
        RECT 25.335 217.320 26.375 217.490 ;
        RECT 26.590 217.460 26.760 217.790 ;
        RECT 27.100 216.920 27.390 218.330 ;
        RECT 24.440 216.880 27.390 216.920 ;
        RECT 17.820 216.680 20.560 216.710 ;
        RECT 14.430 216.290 17.260 216.340 ;
        RECT 14.310 216.170 17.260 216.290 ;
        RECT 14.310 214.760 14.600 216.170 ;
        RECT 14.940 215.300 15.110 215.630 ;
        RECT 15.325 215.600 16.365 215.770 ;
        RECT 15.325 215.160 16.365 215.330 ;
        RECT 16.580 215.300 16.750 215.630 ;
        RECT 17.090 214.760 17.260 216.170 ;
        RECT 14.310 214.640 17.260 214.760 ;
        RECT 14.430 214.590 17.260 214.640 ;
        RECT 17.820 216.260 20.560 216.330 ;
        RECT 21.140 216.320 23.880 216.770 ;
        RECT 17.820 216.160 20.690 216.260 ;
        RECT 17.820 214.750 17.990 216.160 ;
        RECT 18.330 215.290 18.500 215.620 ;
        RECT 18.670 215.590 19.710 215.760 ;
        RECT 18.670 215.150 19.710 215.320 ;
        RECT 19.880 215.290 20.050 215.620 ;
        RECT 20.390 214.750 20.690 216.160 ;
        RECT 17.820 214.610 20.690 214.750 ;
        RECT 21.010 216.220 23.880 216.320 ;
        RECT 24.420 216.800 27.390 216.880 ;
        RECT 24.420 216.350 27.380 216.800 ;
        RECT 24.420 216.270 27.390 216.350 ;
        RECT 21.010 214.810 21.310 216.220 ;
        RECT 21.650 215.350 21.820 215.680 ;
        RECT 21.990 215.650 23.030 215.820 ;
        RECT 21.990 215.210 23.030 215.380 ;
        RECT 23.200 215.350 23.370 215.680 ;
        RECT 23.710 214.810 23.880 216.220 ;
        RECT 21.010 214.670 23.880 214.810 ;
        RECT 17.820 214.580 20.560 214.610 ;
        RECT 14.430 214.190 17.260 214.240 ;
        RECT 14.310 214.070 17.260 214.190 ;
        RECT 14.310 212.660 14.600 214.070 ;
        RECT 14.940 213.200 15.110 213.530 ;
        RECT 15.325 213.500 16.365 213.670 ;
        RECT 15.325 213.060 16.365 213.230 ;
        RECT 16.580 213.200 16.750 213.530 ;
        RECT 17.090 212.660 17.260 214.070 ;
        RECT 14.310 212.540 17.260 212.660 ;
        RECT 14.430 212.490 17.260 212.540 ;
        RECT 17.820 214.160 20.560 214.230 ;
        RECT 21.140 214.220 23.880 214.670 ;
        RECT 24.440 216.230 27.390 216.270 ;
        RECT 24.440 214.820 24.610 216.230 ;
        RECT 24.950 215.360 25.120 215.690 ;
        RECT 25.335 215.660 26.375 215.830 ;
        RECT 25.335 215.220 26.375 215.390 ;
        RECT 26.590 215.360 26.760 215.690 ;
        RECT 27.100 214.820 27.390 216.230 ;
        RECT 24.440 214.700 27.390 214.820 ;
        RECT 24.440 214.650 27.270 214.700 ;
        RECT 17.820 214.060 20.690 214.160 ;
        RECT 17.820 212.650 17.990 214.060 ;
        RECT 18.330 213.190 18.500 213.520 ;
        RECT 18.670 213.490 19.710 213.660 ;
        RECT 18.670 213.050 19.710 213.220 ;
        RECT 19.880 213.190 20.050 213.520 ;
        RECT 20.390 212.650 20.690 214.060 ;
        RECT 17.820 212.510 20.690 212.650 ;
        RECT 21.010 214.120 23.880 214.220 ;
        RECT 21.010 212.710 21.310 214.120 ;
        RECT 21.650 213.250 21.820 213.580 ;
        RECT 21.990 213.550 23.030 213.720 ;
        RECT 21.990 213.110 23.030 213.280 ;
        RECT 23.200 213.250 23.370 213.580 ;
        RECT 23.710 212.710 23.880 214.120 ;
        RECT 21.010 212.570 23.880 212.710 ;
        RECT 21.140 212.540 23.880 212.570 ;
        RECT 24.440 214.250 27.270 214.300 ;
        RECT 24.440 214.130 27.390 214.250 ;
        RECT 24.440 212.720 24.610 214.130 ;
        RECT 24.950 213.260 25.120 213.590 ;
        RECT 25.335 213.560 26.375 213.730 ;
        RECT 25.335 213.120 26.375 213.290 ;
        RECT 26.590 213.260 26.760 213.590 ;
        RECT 27.100 212.720 27.390 214.130 ;
        RECT 24.440 212.600 27.390 212.720 ;
        RECT 24.440 212.550 27.270 212.600 ;
        RECT 17.820 212.480 20.560 212.510 ;
        RECT 14.430 212.100 17.260 212.150 ;
        RECT 14.310 211.980 17.260 212.100 ;
        RECT 14.310 210.570 14.600 211.980 ;
        RECT 14.940 211.110 15.110 211.440 ;
        RECT 15.325 211.410 16.365 211.580 ;
        RECT 15.325 210.970 16.365 211.140 ;
        RECT 16.580 211.110 16.750 211.440 ;
        RECT 17.090 210.570 17.260 211.980 ;
        RECT 14.310 210.450 17.260 210.570 ;
        RECT 14.430 210.400 17.260 210.450 ;
        RECT 17.820 212.070 20.560 212.140 ;
        RECT 21.140 212.120 23.880 212.190 ;
        RECT 17.820 211.970 20.690 212.070 ;
        RECT 17.820 210.560 17.990 211.970 ;
        RECT 18.330 211.100 18.500 211.430 ;
        RECT 18.670 211.400 19.710 211.570 ;
        RECT 18.670 210.960 19.710 211.130 ;
        RECT 19.880 211.100 20.050 211.430 ;
        RECT 20.390 210.560 20.690 211.970 ;
        RECT 17.820 210.420 20.690 210.560 ;
        RECT 21.010 212.020 23.880 212.120 ;
        RECT 21.010 210.610 21.310 212.020 ;
        RECT 21.650 211.150 21.820 211.480 ;
        RECT 21.990 211.450 23.030 211.620 ;
        RECT 21.990 211.010 23.030 211.180 ;
        RECT 23.200 211.150 23.370 211.480 ;
        RECT 23.710 210.610 23.880 212.020 ;
        RECT 21.010 210.470 23.880 210.610 ;
        RECT 21.140 210.440 23.880 210.470 ;
        RECT 24.440 212.150 27.270 212.200 ;
        RECT 24.440 212.030 27.390 212.150 ;
        RECT 24.440 210.620 24.610 212.030 ;
        RECT 24.950 211.160 25.120 211.490 ;
        RECT 25.335 211.460 26.375 211.630 ;
        RECT 25.335 211.020 26.375 211.190 ;
        RECT 26.590 211.160 26.760 211.490 ;
        RECT 27.100 210.620 27.390 212.030 ;
        RECT 24.440 210.500 27.390 210.620 ;
        RECT 24.440 210.450 27.270 210.500 ;
        RECT 17.820 210.390 20.560 210.420 ;
        RECT 14.430 210.000 17.260 210.050 ;
        RECT 14.310 209.880 17.260 210.000 ;
        RECT 14.310 208.470 14.600 209.880 ;
        RECT 14.940 209.010 15.110 209.340 ;
        RECT 15.325 209.310 16.365 209.480 ;
        RECT 15.325 208.870 16.365 209.040 ;
        RECT 16.580 209.010 16.750 209.340 ;
        RECT 17.090 208.470 17.260 209.880 ;
        RECT 14.310 208.350 17.260 208.470 ;
        RECT 14.430 208.300 17.260 208.350 ;
        RECT 17.820 209.970 20.560 210.040 ;
        RECT 21.140 210.020 23.880 210.090 ;
        RECT 17.820 209.870 20.690 209.970 ;
        RECT 17.820 208.460 17.990 209.870 ;
        RECT 18.330 209.000 18.500 209.330 ;
        RECT 18.670 209.300 19.710 209.470 ;
        RECT 18.670 208.860 19.710 209.030 ;
        RECT 19.880 209.000 20.050 209.330 ;
        RECT 20.390 208.460 20.690 209.870 ;
        RECT 17.820 208.320 20.690 208.460 ;
        RECT 21.010 209.920 23.880 210.020 ;
        RECT 21.010 208.510 21.310 209.920 ;
        RECT 21.650 209.050 21.820 209.380 ;
        RECT 21.990 209.350 23.030 209.520 ;
        RECT 21.990 208.910 23.030 209.080 ;
        RECT 23.200 209.050 23.370 209.380 ;
        RECT 23.710 208.510 23.880 209.920 ;
        RECT 21.010 208.370 23.880 208.510 ;
        RECT 21.140 208.340 23.880 208.370 ;
        RECT 24.440 210.050 27.270 210.100 ;
        RECT 24.440 209.930 27.390 210.050 ;
        RECT 24.440 208.520 24.610 209.930 ;
        RECT 24.950 209.060 25.120 209.390 ;
        RECT 25.335 209.360 26.375 209.530 ;
        RECT 25.335 208.920 26.375 209.090 ;
        RECT 26.590 209.060 26.760 209.390 ;
        RECT 27.100 208.520 27.390 209.930 ;
        RECT 24.440 208.400 27.390 208.520 ;
        RECT 24.440 208.350 27.270 208.400 ;
        RECT 17.820 208.290 20.560 208.320 ;
        RECT 14.430 207.910 17.260 207.960 ;
        RECT 14.310 207.790 17.260 207.910 ;
        RECT 14.310 206.380 14.600 207.790 ;
        RECT 14.940 206.920 15.110 207.250 ;
        RECT 15.325 207.220 16.365 207.390 ;
        RECT 15.325 206.780 16.365 206.950 ;
        RECT 16.580 206.920 16.750 207.250 ;
        RECT 17.090 206.380 17.260 207.790 ;
        RECT 14.310 206.260 17.260 206.380 ;
        RECT 14.430 206.210 17.260 206.260 ;
        RECT 17.820 207.880 20.560 207.950 ;
        RECT 21.140 207.920 23.880 207.990 ;
        RECT 17.820 207.780 20.690 207.880 ;
        RECT 17.820 206.370 17.990 207.780 ;
        RECT 18.330 206.910 18.500 207.240 ;
        RECT 18.670 207.210 19.710 207.380 ;
        RECT 18.670 206.770 19.710 206.940 ;
        RECT 19.880 206.910 20.050 207.240 ;
        RECT 20.390 206.370 20.690 207.780 ;
        RECT 17.820 206.230 20.690 206.370 ;
        RECT 21.010 207.820 23.880 207.920 ;
        RECT 21.010 206.410 21.310 207.820 ;
        RECT 21.650 206.950 21.820 207.280 ;
        RECT 21.990 207.250 23.030 207.420 ;
        RECT 21.990 206.810 23.030 206.980 ;
        RECT 23.200 206.950 23.370 207.280 ;
        RECT 23.710 206.410 23.880 207.820 ;
        RECT 21.010 206.270 23.880 206.410 ;
        RECT 21.140 206.240 23.880 206.270 ;
        RECT 24.440 207.950 27.270 208.000 ;
        RECT 24.440 207.830 27.390 207.950 ;
        RECT 24.440 206.420 24.610 207.830 ;
        RECT 24.950 206.960 25.120 207.290 ;
        RECT 25.335 207.260 26.375 207.430 ;
        RECT 25.335 206.820 26.375 206.990 ;
        RECT 26.590 206.960 26.760 207.290 ;
        RECT 27.100 206.420 27.390 207.830 ;
        RECT 24.440 206.300 27.390 206.420 ;
        RECT 24.440 206.250 27.270 206.300 ;
        RECT 17.820 206.200 20.560 206.230 ;
        RECT 14.430 205.810 17.260 205.860 ;
        RECT 14.310 205.690 17.260 205.810 ;
        RECT 14.310 204.280 14.600 205.690 ;
        RECT 14.940 204.820 15.110 205.150 ;
        RECT 15.325 205.120 16.365 205.290 ;
        RECT 15.325 204.680 16.365 204.850 ;
        RECT 16.580 204.820 16.750 205.150 ;
        RECT 17.090 204.280 17.260 205.690 ;
        RECT 14.310 204.160 17.260 204.280 ;
        RECT 14.430 204.110 17.260 204.160 ;
        RECT 17.820 205.780 20.560 205.850 ;
        RECT 21.140 205.820 23.880 205.890 ;
        RECT 17.820 205.680 20.690 205.780 ;
        RECT 17.820 204.270 17.990 205.680 ;
        RECT 18.330 204.810 18.500 205.140 ;
        RECT 18.670 205.110 19.710 205.280 ;
        RECT 18.670 204.670 19.710 204.840 ;
        RECT 19.880 204.810 20.050 205.140 ;
        RECT 20.390 204.270 20.690 205.680 ;
        RECT 17.820 204.130 20.690 204.270 ;
        RECT 21.010 205.720 23.880 205.820 ;
        RECT 21.010 204.310 21.310 205.720 ;
        RECT 21.650 204.850 21.820 205.180 ;
        RECT 21.990 205.150 23.030 205.320 ;
        RECT 21.990 204.710 23.030 204.880 ;
        RECT 23.200 204.850 23.370 205.180 ;
        RECT 23.710 204.310 23.880 205.720 ;
        RECT 21.010 204.170 23.880 204.310 ;
        RECT 21.140 204.140 23.880 204.170 ;
        RECT 24.440 205.850 27.270 205.900 ;
        RECT 24.440 205.730 27.390 205.850 ;
        RECT 24.440 204.320 24.610 205.730 ;
        RECT 24.950 204.860 25.120 205.190 ;
        RECT 25.335 205.160 26.375 205.330 ;
        RECT 25.335 204.720 26.375 204.890 ;
        RECT 26.590 204.860 26.760 205.190 ;
        RECT 27.100 204.320 27.390 205.730 ;
        RECT 24.440 204.200 27.390 204.320 ;
        RECT 24.440 204.150 27.270 204.200 ;
        RECT 17.820 204.100 20.560 204.130 ;
        RECT 14.430 203.710 17.260 203.760 ;
        RECT 14.310 203.590 17.260 203.710 ;
        RECT 14.310 202.180 14.600 203.590 ;
        RECT 14.940 202.720 15.110 203.050 ;
        RECT 15.325 203.020 16.365 203.190 ;
        RECT 15.325 202.580 16.365 202.750 ;
        RECT 16.580 202.720 16.750 203.050 ;
        RECT 17.090 202.180 17.260 203.590 ;
        RECT 14.310 202.060 17.260 202.180 ;
        RECT 14.430 202.010 17.260 202.060 ;
        RECT 17.820 203.680 20.560 203.750 ;
        RECT 21.140 203.720 23.880 203.790 ;
        RECT 17.820 203.580 20.690 203.680 ;
        RECT 17.820 202.170 17.990 203.580 ;
        RECT 18.330 202.710 18.500 203.040 ;
        RECT 18.670 203.010 19.710 203.180 ;
        RECT 18.670 202.570 19.710 202.740 ;
        RECT 19.880 202.710 20.050 203.040 ;
        RECT 20.390 202.170 20.690 203.580 ;
        RECT 17.820 202.030 20.690 202.170 ;
        RECT 21.010 203.620 23.880 203.720 ;
        RECT 21.010 202.210 21.310 203.620 ;
        RECT 21.650 202.750 21.820 203.080 ;
        RECT 21.990 203.050 23.030 203.220 ;
        RECT 21.990 202.610 23.030 202.780 ;
        RECT 23.200 202.750 23.370 203.080 ;
        RECT 23.710 202.210 23.880 203.620 ;
        RECT 21.010 202.070 23.880 202.210 ;
        RECT 21.140 202.040 23.880 202.070 ;
        RECT 24.440 203.750 27.270 203.800 ;
        RECT 24.440 203.630 27.390 203.750 ;
        RECT 24.440 202.220 24.610 203.630 ;
        RECT 24.950 202.760 25.120 203.090 ;
        RECT 25.335 203.060 26.375 203.230 ;
        RECT 25.335 202.620 26.375 202.790 ;
        RECT 26.590 202.760 26.760 203.090 ;
        RECT 27.100 202.220 27.390 203.630 ;
        RECT 24.440 202.100 27.390 202.220 ;
        RECT 24.440 202.050 27.270 202.100 ;
        RECT 17.820 202.000 20.560 202.030 ;
        RECT 14.430 201.610 17.260 201.660 ;
        RECT 14.310 201.490 17.260 201.610 ;
        RECT 14.310 200.080 14.600 201.490 ;
        RECT 14.940 200.620 15.110 200.950 ;
        RECT 15.325 200.920 16.365 201.090 ;
        RECT 15.325 200.480 16.365 200.650 ;
        RECT 16.580 200.620 16.750 200.950 ;
        RECT 17.090 200.080 17.260 201.490 ;
        RECT 14.310 199.960 17.260 200.080 ;
        RECT 14.430 199.910 17.260 199.960 ;
        RECT 17.820 201.580 20.560 201.650 ;
        RECT 21.140 201.620 23.880 201.690 ;
        RECT 17.820 201.480 20.690 201.580 ;
        RECT 17.820 200.070 17.990 201.480 ;
        RECT 18.330 200.610 18.500 200.940 ;
        RECT 18.670 200.910 19.710 201.080 ;
        RECT 18.670 200.470 19.710 200.640 ;
        RECT 19.880 200.610 20.050 200.940 ;
        RECT 20.390 200.070 20.690 201.480 ;
        RECT 17.820 199.930 20.690 200.070 ;
        RECT 21.010 201.520 23.880 201.620 ;
        RECT 21.010 200.110 21.310 201.520 ;
        RECT 21.650 200.650 21.820 200.980 ;
        RECT 21.990 200.950 23.030 201.120 ;
        RECT 21.990 200.510 23.030 200.680 ;
        RECT 23.200 200.650 23.370 200.980 ;
        RECT 23.710 200.110 23.880 201.520 ;
        RECT 21.010 199.970 23.880 200.110 ;
        RECT 21.140 199.940 23.880 199.970 ;
        RECT 24.440 201.650 27.270 201.700 ;
        RECT 24.440 201.530 27.390 201.650 ;
        RECT 24.440 200.120 24.610 201.530 ;
        RECT 24.950 200.660 25.120 200.990 ;
        RECT 25.335 200.960 26.375 201.130 ;
        RECT 25.335 200.520 26.375 200.690 ;
        RECT 26.590 200.660 26.760 200.990 ;
        RECT 27.100 200.120 27.390 201.530 ;
        RECT 24.440 200.000 27.390 200.120 ;
        RECT 24.440 199.950 27.270 200.000 ;
        RECT 17.820 199.900 20.560 199.930 ;
        RECT 14.430 199.510 17.260 199.560 ;
        RECT 14.310 199.390 17.260 199.510 ;
        RECT 14.310 197.980 14.600 199.390 ;
        RECT 14.940 198.520 15.110 198.850 ;
        RECT 15.325 198.820 16.365 198.990 ;
        RECT 15.325 198.380 16.365 198.550 ;
        RECT 16.580 198.520 16.750 198.850 ;
        RECT 17.090 197.980 17.260 199.390 ;
        RECT 14.310 197.860 17.260 197.980 ;
        RECT 14.430 197.810 17.260 197.860 ;
        RECT 17.820 199.480 20.560 199.550 ;
        RECT 21.140 199.520 23.880 199.590 ;
        RECT 17.820 199.380 20.690 199.480 ;
        RECT 17.820 197.970 17.990 199.380 ;
        RECT 18.330 198.510 18.500 198.840 ;
        RECT 18.670 198.810 19.710 198.980 ;
        RECT 18.670 198.370 19.710 198.540 ;
        RECT 19.880 198.510 20.050 198.840 ;
        RECT 20.390 197.970 20.690 199.380 ;
        RECT 17.820 197.830 20.690 197.970 ;
        RECT 21.010 199.420 23.880 199.520 ;
        RECT 21.010 198.010 21.310 199.420 ;
        RECT 21.650 198.550 21.820 198.880 ;
        RECT 21.990 198.850 23.030 199.020 ;
        RECT 21.990 198.410 23.030 198.580 ;
        RECT 23.200 198.550 23.370 198.880 ;
        RECT 23.710 198.010 23.880 199.420 ;
        RECT 21.010 197.870 23.880 198.010 ;
        RECT 21.140 197.840 23.880 197.870 ;
        RECT 24.440 199.550 27.270 199.600 ;
        RECT 24.440 199.430 27.390 199.550 ;
        RECT 24.440 198.020 24.610 199.430 ;
        RECT 24.950 198.560 25.120 198.890 ;
        RECT 25.335 198.860 26.375 199.030 ;
        RECT 25.335 198.420 26.375 198.590 ;
        RECT 26.590 198.560 26.760 198.890 ;
        RECT 27.100 198.020 27.390 199.430 ;
        RECT 24.440 197.900 27.390 198.020 ;
        RECT 24.440 197.850 27.270 197.900 ;
        RECT 17.820 197.800 20.560 197.830 ;
        RECT 14.430 197.410 17.260 197.460 ;
        RECT 14.310 197.290 17.260 197.410 ;
        RECT 14.310 195.880 14.600 197.290 ;
        RECT 14.940 196.420 15.110 196.750 ;
        RECT 15.325 196.720 16.365 196.890 ;
        RECT 15.325 196.280 16.365 196.450 ;
        RECT 16.580 196.420 16.750 196.750 ;
        RECT 17.090 195.880 17.260 197.290 ;
        RECT 14.310 195.760 17.260 195.880 ;
        RECT 14.430 195.710 17.260 195.760 ;
        RECT 17.820 197.380 20.560 197.450 ;
        RECT 21.140 197.420 23.880 197.490 ;
        RECT 17.820 197.280 20.690 197.380 ;
        RECT 17.820 195.870 17.990 197.280 ;
        RECT 18.330 196.410 18.500 196.740 ;
        RECT 18.670 196.710 19.710 196.880 ;
        RECT 18.670 196.270 19.710 196.440 ;
        RECT 19.880 196.410 20.050 196.740 ;
        RECT 20.390 195.870 20.690 197.280 ;
        RECT 17.820 195.730 20.690 195.870 ;
        RECT 21.010 197.320 23.880 197.420 ;
        RECT 21.010 195.910 21.310 197.320 ;
        RECT 21.650 196.450 21.820 196.780 ;
        RECT 21.990 196.750 23.030 196.920 ;
        RECT 21.990 196.310 23.030 196.480 ;
        RECT 23.200 196.450 23.370 196.780 ;
        RECT 23.710 195.910 23.880 197.320 ;
        RECT 21.010 195.770 23.880 195.910 ;
        RECT 21.140 195.740 23.880 195.770 ;
        RECT 24.440 197.450 27.270 197.500 ;
        RECT 24.440 197.330 27.390 197.450 ;
        RECT 24.440 195.920 24.610 197.330 ;
        RECT 24.950 196.460 25.120 196.790 ;
        RECT 25.335 196.760 26.375 196.930 ;
        RECT 25.335 196.320 26.375 196.490 ;
        RECT 26.590 196.460 26.760 196.790 ;
        RECT 27.100 195.920 27.390 197.330 ;
        RECT 24.440 195.800 27.390 195.920 ;
        RECT 24.440 195.750 27.270 195.800 ;
        RECT 17.820 195.700 20.560 195.730 ;
        RECT 14.430 195.310 17.260 195.360 ;
        RECT 14.310 195.190 17.260 195.310 ;
        RECT 14.310 193.780 14.600 195.190 ;
        RECT 14.940 194.320 15.110 194.650 ;
        RECT 15.325 194.620 16.365 194.790 ;
        RECT 15.325 194.180 16.365 194.350 ;
        RECT 16.580 194.320 16.750 194.650 ;
        RECT 17.090 193.780 17.260 195.190 ;
        RECT 14.310 193.660 17.260 193.780 ;
        RECT 14.430 193.610 17.260 193.660 ;
        RECT 17.820 195.280 20.560 195.350 ;
        RECT 21.140 195.320 23.880 195.390 ;
        RECT 17.820 195.180 20.690 195.280 ;
        RECT 17.820 193.770 17.990 195.180 ;
        RECT 18.330 194.310 18.500 194.640 ;
        RECT 18.670 194.610 19.710 194.780 ;
        RECT 18.670 194.170 19.710 194.340 ;
        RECT 19.880 194.310 20.050 194.640 ;
        RECT 20.390 193.770 20.690 195.180 ;
        RECT 17.820 193.630 20.690 193.770 ;
        RECT 21.010 195.220 23.880 195.320 ;
        RECT 21.010 193.810 21.310 195.220 ;
        RECT 21.650 194.350 21.820 194.680 ;
        RECT 21.990 194.650 23.030 194.820 ;
        RECT 21.990 194.210 23.030 194.380 ;
        RECT 23.200 194.350 23.370 194.680 ;
        RECT 23.710 193.810 23.880 195.220 ;
        RECT 21.010 193.670 23.880 193.810 ;
        RECT 21.140 193.640 23.880 193.670 ;
        RECT 24.440 195.350 27.270 195.400 ;
        RECT 24.440 195.230 27.390 195.350 ;
        RECT 24.440 193.820 24.610 195.230 ;
        RECT 24.950 194.360 25.120 194.690 ;
        RECT 25.335 194.660 26.375 194.830 ;
        RECT 25.335 194.220 26.375 194.390 ;
        RECT 26.590 194.360 26.760 194.690 ;
        RECT 27.100 193.820 27.390 195.230 ;
        RECT 24.440 193.700 27.390 193.820 ;
        RECT 24.440 193.650 27.270 193.700 ;
        RECT 17.820 193.600 20.560 193.630 ;
        RECT 14.430 193.210 17.260 193.260 ;
        RECT 14.310 193.090 17.260 193.210 ;
        RECT 14.310 191.680 14.600 193.090 ;
        RECT 14.940 192.220 15.110 192.550 ;
        RECT 15.325 192.520 16.365 192.690 ;
        RECT 15.325 192.080 16.365 192.250 ;
        RECT 16.580 192.220 16.750 192.550 ;
        RECT 17.090 191.680 17.260 193.090 ;
        RECT 14.310 191.560 17.260 191.680 ;
        RECT 14.430 191.510 17.260 191.560 ;
        RECT 17.820 193.180 20.560 193.250 ;
        RECT 21.140 193.220 23.880 193.290 ;
        RECT 17.820 193.080 20.690 193.180 ;
        RECT 17.820 191.670 17.990 193.080 ;
        RECT 18.330 192.210 18.500 192.540 ;
        RECT 18.670 192.510 19.710 192.680 ;
        RECT 18.670 192.070 19.710 192.240 ;
        RECT 19.880 192.210 20.050 192.540 ;
        RECT 20.390 191.670 20.690 193.080 ;
        RECT 17.820 191.530 20.690 191.670 ;
        RECT 21.010 193.120 23.880 193.220 ;
        RECT 21.010 191.710 21.310 193.120 ;
        RECT 21.650 192.250 21.820 192.580 ;
        RECT 21.990 192.550 23.030 192.720 ;
        RECT 21.990 192.110 23.030 192.280 ;
        RECT 23.200 192.250 23.370 192.580 ;
        RECT 23.710 191.710 23.880 193.120 ;
        RECT 21.010 191.570 23.880 191.710 ;
        RECT 21.140 191.540 23.880 191.570 ;
        RECT 24.440 193.250 27.270 193.300 ;
        RECT 24.440 193.130 27.390 193.250 ;
        RECT 24.440 191.720 24.610 193.130 ;
        RECT 24.950 192.260 25.120 192.590 ;
        RECT 25.335 192.560 26.375 192.730 ;
        RECT 25.335 192.120 26.375 192.290 ;
        RECT 26.590 192.260 26.760 192.590 ;
        RECT 27.100 191.720 27.390 193.130 ;
        RECT 24.440 191.600 27.390 191.720 ;
        RECT 24.440 191.550 27.270 191.600 ;
        RECT 17.820 191.500 20.560 191.530 ;
        RECT 14.430 191.110 17.260 191.160 ;
        RECT 14.310 190.990 17.260 191.110 ;
        RECT 14.310 189.580 14.600 190.990 ;
        RECT 14.940 190.120 15.110 190.450 ;
        RECT 15.325 190.420 16.365 190.590 ;
        RECT 15.325 189.980 16.365 190.150 ;
        RECT 16.580 190.120 16.750 190.450 ;
        RECT 17.090 189.580 17.260 190.990 ;
        RECT 14.310 189.460 17.260 189.580 ;
        RECT 14.430 189.410 17.260 189.460 ;
        RECT 17.820 191.080 20.560 191.150 ;
        RECT 21.140 191.120 23.880 191.190 ;
        RECT 17.820 190.980 20.690 191.080 ;
        RECT 17.820 189.570 17.990 190.980 ;
        RECT 18.330 190.110 18.500 190.440 ;
        RECT 18.670 190.410 19.710 190.580 ;
        RECT 18.670 189.970 19.710 190.140 ;
        RECT 19.880 190.110 20.050 190.440 ;
        RECT 20.390 189.570 20.690 190.980 ;
        RECT 17.820 189.430 20.690 189.570 ;
        RECT 21.010 191.020 23.880 191.120 ;
        RECT 21.010 189.610 21.310 191.020 ;
        RECT 21.650 190.150 21.820 190.480 ;
        RECT 21.990 190.450 23.030 190.620 ;
        RECT 21.990 190.010 23.030 190.180 ;
        RECT 23.200 190.150 23.370 190.480 ;
        RECT 23.710 189.610 23.880 191.020 ;
        RECT 21.010 189.470 23.880 189.610 ;
        RECT 21.140 189.440 23.880 189.470 ;
        RECT 24.440 191.150 27.270 191.200 ;
        RECT 24.440 191.030 27.390 191.150 ;
        RECT 24.440 189.620 24.610 191.030 ;
        RECT 24.950 190.160 25.120 190.490 ;
        RECT 25.335 190.460 26.375 190.630 ;
        RECT 25.335 190.020 26.375 190.190 ;
        RECT 26.590 190.160 26.760 190.490 ;
        RECT 27.100 189.620 27.390 191.030 ;
        RECT 24.440 189.500 27.390 189.620 ;
        RECT 24.440 189.450 27.270 189.500 ;
        RECT 17.820 189.400 20.560 189.430 ;
        RECT 14.430 189.020 17.260 189.070 ;
        RECT 14.310 188.900 17.260 189.020 ;
        RECT 14.310 187.490 14.600 188.900 ;
        RECT 14.940 188.030 15.110 188.360 ;
        RECT 15.325 188.330 16.365 188.500 ;
        RECT 15.325 187.890 16.365 188.060 ;
        RECT 16.580 188.030 16.750 188.360 ;
        RECT 17.090 187.490 17.260 188.900 ;
        RECT 14.310 187.370 17.260 187.490 ;
        RECT 14.430 187.320 17.260 187.370 ;
        RECT 17.820 188.990 20.560 189.060 ;
        RECT 21.140 189.020 23.880 189.090 ;
        RECT 17.820 188.890 20.690 188.990 ;
        RECT 17.820 187.480 17.990 188.890 ;
        RECT 18.330 188.020 18.500 188.350 ;
        RECT 18.670 188.320 19.710 188.490 ;
        RECT 18.670 187.880 19.710 188.050 ;
        RECT 19.880 188.020 20.050 188.350 ;
        RECT 20.390 187.480 20.690 188.890 ;
        RECT 17.820 187.340 20.690 187.480 ;
        RECT 21.010 188.920 23.880 189.020 ;
        RECT 21.010 187.510 21.310 188.920 ;
        RECT 21.650 188.050 21.820 188.380 ;
        RECT 21.990 188.350 23.030 188.520 ;
        RECT 21.990 187.910 23.030 188.080 ;
        RECT 23.200 188.050 23.370 188.380 ;
        RECT 23.710 187.510 23.880 188.920 ;
        RECT 21.010 187.370 23.880 187.510 ;
        RECT 21.140 187.340 23.880 187.370 ;
        RECT 24.440 189.050 27.270 189.100 ;
        RECT 24.440 188.930 27.390 189.050 ;
        RECT 24.440 187.520 24.610 188.930 ;
        RECT 24.950 188.060 25.120 188.390 ;
        RECT 25.335 188.360 26.375 188.530 ;
        RECT 25.335 187.920 26.375 188.090 ;
        RECT 26.590 188.060 26.760 188.390 ;
        RECT 27.100 187.520 27.390 188.930 ;
        RECT 24.440 187.400 27.390 187.520 ;
        RECT 24.440 187.350 27.270 187.400 ;
        RECT 17.820 187.310 20.560 187.340 ;
        RECT 14.430 186.930 17.260 186.980 ;
        RECT 14.310 186.810 17.260 186.930 ;
        RECT 14.310 185.400 14.600 186.810 ;
        RECT 14.940 185.940 15.110 186.270 ;
        RECT 15.325 186.240 16.365 186.410 ;
        RECT 15.325 185.800 16.365 185.970 ;
        RECT 16.580 185.940 16.750 186.270 ;
        RECT 17.090 185.400 17.260 186.810 ;
        RECT 14.310 185.280 17.260 185.400 ;
        RECT 14.430 185.230 17.260 185.280 ;
        RECT 17.820 186.900 20.560 186.970 ;
        RECT 21.140 186.920 23.880 186.990 ;
        RECT 17.820 186.800 20.690 186.900 ;
        RECT 17.820 185.390 17.990 186.800 ;
        RECT 18.330 185.930 18.500 186.260 ;
        RECT 18.670 186.230 19.710 186.400 ;
        RECT 18.670 185.790 19.710 185.960 ;
        RECT 19.880 185.930 20.050 186.260 ;
        RECT 20.390 185.390 20.690 186.800 ;
        RECT 17.820 185.250 20.690 185.390 ;
        RECT 21.010 186.820 23.880 186.920 ;
        RECT 21.010 185.410 21.310 186.820 ;
        RECT 21.650 185.950 21.820 186.280 ;
        RECT 21.990 186.250 23.030 186.420 ;
        RECT 21.990 185.810 23.030 185.980 ;
        RECT 23.200 185.950 23.370 186.280 ;
        RECT 23.710 185.410 23.880 186.820 ;
        RECT 21.010 185.270 23.880 185.410 ;
        RECT 17.820 185.220 20.560 185.250 ;
        RECT 21.140 185.240 23.880 185.270 ;
        RECT 24.440 186.950 27.270 187.000 ;
        RECT 24.440 186.830 27.390 186.950 ;
        RECT 24.440 185.420 24.610 186.830 ;
        RECT 24.950 185.960 25.120 186.290 ;
        RECT 25.335 186.260 26.375 186.430 ;
        RECT 25.335 185.820 26.375 185.990 ;
        RECT 26.590 185.960 26.760 186.290 ;
        RECT 27.100 185.420 27.390 186.830 ;
        RECT 24.440 185.300 27.390 185.420 ;
        RECT 24.440 185.250 27.270 185.300 ;
        RECT 14.430 184.830 17.260 184.880 ;
        RECT 14.310 184.710 17.260 184.830 ;
        RECT 14.310 183.300 14.600 184.710 ;
        RECT 14.940 183.840 15.110 184.170 ;
        RECT 15.325 184.140 16.365 184.310 ;
        RECT 15.325 183.700 16.365 183.870 ;
        RECT 16.580 183.840 16.750 184.170 ;
        RECT 17.090 183.300 17.260 184.710 ;
        RECT 14.310 183.180 17.260 183.300 ;
        RECT 14.430 183.130 17.260 183.180 ;
        RECT 17.820 184.800 20.560 184.870 ;
        RECT 21.140 184.820 23.880 184.890 ;
        RECT 17.820 184.700 20.690 184.800 ;
        RECT 17.820 183.290 17.990 184.700 ;
        RECT 18.330 183.830 18.500 184.160 ;
        RECT 18.670 184.130 19.710 184.300 ;
        RECT 18.670 183.690 19.710 183.860 ;
        RECT 19.880 183.830 20.050 184.160 ;
        RECT 20.390 183.290 20.690 184.700 ;
        RECT 17.820 183.150 20.690 183.290 ;
        RECT 21.010 184.720 23.880 184.820 ;
        RECT 21.010 183.310 21.310 184.720 ;
        RECT 21.650 183.850 21.820 184.180 ;
        RECT 21.990 184.150 23.030 184.320 ;
        RECT 21.990 183.710 23.030 183.880 ;
        RECT 23.200 183.850 23.370 184.180 ;
        RECT 23.710 183.310 23.880 184.720 ;
        RECT 21.010 183.170 23.880 183.310 ;
        RECT 17.820 183.120 20.560 183.150 ;
        RECT 21.140 183.140 23.880 183.170 ;
        RECT 24.440 184.850 27.270 184.900 ;
        RECT 24.440 184.730 27.390 184.850 ;
        RECT 24.440 183.320 24.610 184.730 ;
        RECT 24.950 183.860 25.120 184.190 ;
        RECT 25.335 184.160 26.375 184.330 ;
        RECT 25.335 183.720 26.375 183.890 ;
        RECT 26.590 183.860 26.760 184.190 ;
        RECT 27.100 183.320 27.390 184.730 ;
        RECT 24.440 183.200 27.390 183.320 ;
        RECT 24.440 183.150 27.270 183.200 ;
        RECT 14.430 182.740 17.260 182.790 ;
        RECT 14.310 182.620 17.260 182.740 ;
        RECT 14.310 181.210 14.600 182.620 ;
        RECT 14.940 181.750 15.110 182.080 ;
        RECT 15.325 182.050 16.365 182.220 ;
        RECT 15.325 181.610 16.365 181.780 ;
        RECT 16.580 181.750 16.750 182.080 ;
        RECT 17.090 181.210 17.260 182.620 ;
        RECT 14.310 181.090 17.260 181.210 ;
        RECT 14.430 181.040 17.260 181.090 ;
        RECT 17.820 182.710 20.560 182.780 ;
        RECT 21.140 182.720 23.880 182.790 ;
        RECT 17.820 182.610 20.690 182.710 ;
        RECT 17.820 181.200 17.990 182.610 ;
        RECT 18.330 181.740 18.500 182.070 ;
        RECT 18.670 182.040 19.710 182.210 ;
        RECT 18.670 181.600 19.710 181.770 ;
        RECT 19.880 181.740 20.050 182.070 ;
        RECT 20.390 181.200 20.690 182.610 ;
        RECT 17.820 181.060 20.690 181.200 ;
        RECT 21.010 182.620 23.880 182.720 ;
        RECT 21.010 181.210 21.310 182.620 ;
        RECT 21.650 181.750 21.820 182.080 ;
        RECT 21.990 182.050 23.030 182.220 ;
        RECT 21.990 181.610 23.030 181.780 ;
        RECT 23.200 181.750 23.370 182.080 ;
        RECT 23.710 181.210 23.880 182.620 ;
        RECT 21.010 181.070 23.880 181.210 ;
        RECT 17.820 181.030 20.560 181.060 ;
        RECT 21.140 181.040 23.880 181.070 ;
        RECT 24.440 182.750 27.270 182.800 ;
        RECT 24.440 182.630 27.390 182.750 ;
        RECT 24.440 181.220 24.610 182.630 ;
        RECT 24.950 181.760 25.120 182.090 ;
        RECT 25.335 182.060 26.375 182.230 ;
        RECT 25.335 181.620 26.375 181.790 ;
        RECT 26.590 181.760 26.760 182.090 ;
        RECT 27.100 181.220 27.390 182.630 ;
        RECT 24.440 181.100 27.390 181.220 ;
        RECT 24.440 181.050 27.270 181.100 ;
        RECT 14.430 180.650 17.260 180.700 ;
        RECT 14.310 180.530 17.260 180.650 ;
        RECT 14.310 179.120 14.600 180.530 ;
        RECT 14.940 179.660 15.110 179.990 ;
        RECT 15.325 179.960 16.365 180.130 ;
        RECT 15.325 179.520 16.365 179.690 ;
        RECT 16.580 179.660 16.750 179.990 ;
        RECT 17.090 179.120 17.260 180.530 ;
        RECT 14.310 179.000 17.260 179.120 ;
        RECT 14.430 178.950 17.260 179.000 ;
        RECT 17.820 180.620 20.560 180.690 ;
        RECT 21.140 180.620 23.880 180.690 ;
        RECT 17.820 180.520 20.690 180.620 ;
        RECT 17.820 179.110 17.990 180.520 ;
        RECT 18.330 179.650 18.500 179.980 ;
        RECT 18.670 179.950 19.710 180.120 ;
        RECT 18.670 179.510 19.710 179.680 ;
        RECT 19.880 179.650 20.050 179.980 ;
        RECT 20.390 179.110 20.690 180.520 ;
        RECT 17.820 178.970 20.690 179.110 ;
        RECT 21.010 180.520 23.880 180.620 ;
        RECT 21.010 179.110 21.310 180.520 ;
        RECT 21.650 179.650 21.820 179.980 ;
        RECT 21.990 179.950 23.030 180.120 ;
        RECT 21.990 179.510 23.030 179.680 ;
        RECT 23.200 179.650 23.370 179.980 ;
        RECT 23.710 179.110 23.880 180.520 ;
        RECT 21.010 178.970 23.880 179.110 ;
        RECT 17.820 178.940 20.560 178.970 ;
        RECT 21.140 178.940 23.880 178.970 ;
        RECT 24.440 180.650 27.270 180.700 ;
        RECT 24.440 180.530 27.390 180.650 ;
        RECT 24.440 179.120 24.610 180.530 ;
        RECT 24.950 179.660 25.120 179.990 ;
        RECT 25.335 179.960 26.375 180.130 ;
        RECT 25.335 179.520 26.375 179.690 ;
        RECT 26.590 179.660 26.760 179.990 ;
        RECT 27.100 179.120 27.390 180.530 ;
        RECT 24.440 179.000 27.390 179.120 ;
        RECT 24.440 178.950 27.270 179.000 ;
        RECT 14.430 178.550 17.260 178.600 ;
        RECT 14.310 178.430 17.260 178.550 ;
        RECT 14.310 177.020 14.600 178.430 ;
        RECT 14.940 177.560 15.110 177.890 ;
        RECT 15.325 177.860 16.365 178.030 ;
        RECT 15.325 177.420 16.365 177.590 ;
        RECT 16.580 177.560 16.750 177.890 ;
        RECT 17.090 177.020 17.260 178.430 ;
        RECT 14.310 176.900 17.260 177.020 ;
        RECT 14.430 176.850 17.260 176.900 ;
        RECT 17.820 178.520 20.560 178.590 ;
        RECT 21.140 178.520 23.880 178.590 ;
        RECT 17.820 178.420 20.690 178.520 ;
        RECT 17.820 177.010 17.990 178.420 ;
        RECT 18.330 177.550 18.500 177.880 ;
        RECT 18.670 177.850 19.710 178.020 ;
        RECT 18.670 177.410 19.710 177.580 ;
        RECT 19.880 177.550 20.050 177.880 ;
        RECT 20.390 177.010 20.690 178.420 ;
        RECT 17.820 176.870 20.690 177.010 ;
        RECT 21.010 178.420 23.880 178.520 ;
        RECT 21.010 177.010 21.310 178.420 ;
        RECT 21.650 177.550 21.820 177.880 ;
        RECT 21.990 177.850 23.030 178.020 ;
        RECT 21.990 177.410 23.030 177.580 ;
        RECT 23.200 177.550 23.370 177.880 ;
        RECT 23.710 177.010 23.880 178.420 ;
        RECT 21.010 176.870 23.880 177.010 ;
        RECT 17.820 176.840 20.560 176.870 ;
        RECT 21.140 176.840 23.880 176.870 ;
        RECT 24.440 178.550 27.270 178.600 ;
        RECT 24.440 178.430 27.390 178.550 ;
        RECT 24.440 177.020 24.610 178.430 ;
        RECT 24.950 177.560 25.120 177.890 ;
        RECT 25.335 177.860 26.375 178.030 ;
        RECT 25.335 177.420 26.375 177.590 ;
        RECT 26.590 177.560 26.760 177.890 ;
        RECT 27.100 177.020 27.390 178.430 ;
        RECT 24.440 176.900 27.390 177.020 ;
        RECT 24.440 176.850 27.270 176.900 ;
        RECT 14.430 176.450 17.260 176.500 ;
        RECT 14.310 176.330 17.260 176.450 ;
        RECT 14.310 174.920 14.600 176.330 ;
        RECT 14.940 175.460 15.110 175.790 ;
        RECT 15.325 175.760 16.365 175.930 ;
        RECT 15.325 175.320 16.365 175.490 ;
        RECT 16.580 175.460 16.750 175.790 ;
        RECT 17.090 174.920 17.260 176.330 ;
        RECT 14.310 174.800 17.260 174.920 ;
        RECT 14.430 174.750 17.260 174.800 ;
        RECT 17.820 176.420 20.560 176.490 ;
        RECT 21.140 176.420 23.880 176.490 ;
        RECT 17.820 176.320 20.690 176.420 ;
        RECT 17.820 174.910 17.990 176.320 ;
        RECT 18.330 175.450 18.500 175.780 ;
        RECT 18.670 175.750 19.710 175.920 ;
        RECT 18.670 175.310 19.710 175.480 ;
        RECT 19.880 175.450 20.050 175.780 ;
        RECT 20.390 174.910 20.690 176.320 ;
        RECT 17.820 174.770 20.690 174.910 ;
        RECT 21.010 176.320 23.880 176.420 ;
        RECT 21.010 174.910 21.310 176.320 ;
        RECT 21.650 175.450 21.820 175.780 ;
        RECT 21.990 175.750 23.030 175.920 ;
        RECT 21.990 175.310 23.030 175.480 ;
        RECT 23.200 175.450 23.370 175.780 ;
        RECT 23.710 174.910 23.880 176.320 ;
        RECT 21.010 174.770 23.880 174.910 ;
        RECT 17.820 174.740 20.560 174.770 ;
        RECT 21.140 174.740 23.880 174.770 ;
        RECT 24.440 176.450 27.270 176.500 ;
        RECT 24.440 176.330 27.390 176.450 ;
        RECT 24.440 174.920 24.610 176.330 ;
        RECT 24.950 175.460 25.120 175.790 ;
        RECT 25.335 175.760 26.375 175.930 ;
        RECT 25.335 175.320 26.375 175.490 ;
        RECT 26.590 175.460 26.760 175.790 ;
        RECT 27.100 174.920 27.390 176.330 ;
        RECT 24.440 174.800 27.390 174.920 ;
        RECT 24.440 174.750 27.270 174.800 ;
        RECT 14.430 174.350 17.260 174.400 ;
        RECT 14.310 174.230 17.260 174.350 ;
        RECT 14.310 172.820 14.600 174.230 ;
        RECT 14.940 173.360 15.110 173.690 ;
        RECT 15.325 173.660 16.365 173.830 ;
        RECT 15.325 173.220 16.365 173.390 ;
        RECT 16.580 173.360 16.750 173.690 ;
        RECT 17.090 172.820 17.260 174.230 ;
        RECT 14.310 172.700 17.260 172.820 ;
        RECT 14.430 172.650 17.260 172.700 ;
        RECT 17.820 174.320 20.560 174.390 ;
        RECT 21.140 174.320 23.880 174.390 ;
        RECT 17.820 174.220 20.690 174.320 ;
        RECT 17.820 172.810 17.990 174.220 ;
        RECT 18.330 173.350 18.500 173.680 ;
        RECT 18.670 173.650 19.710 173.820 ;
        RECT 18.670 173.210 19.710 173.380 ;
        RECT 19.880 173.350 20.050 173.680 ;
        RECT 20.390 172.810 20.690 174.220 ;
        RECT 17.820 172.670 20.690 172.810 ;
        RECT 21.010 174.220 23.880 174.320 ;
        RECT 21.010 172.810 21.310 174.220 ;
        RECT 21.650 173.350 21.820 173.680 ;
        RECT 21.990 173.650 23.030 173.820 ;
        RECT 21.990 173.210 23.030 173.380 ;
        RECT 23.200 173.350 23.370 173.680 ;
        RECT 23.710 172.810 23.880 174.220 ;
        RECT 21.010 172.670 23.880 172.810 ;
        RECT 17.820 172.640 20.560 172.670 ;
        RECT 21.140 172.640 23.880 172.670 ;
        RECT 24.440 174.350 27.270 174.400 ;
        RECT 24.440 174.230 27.390 174.350 ;
        RECT 24.440 172.820 24.610 174.230 ;
        RECT 24.950 173.360 25.120 173.690 ;
        RECT 25.335 173.660 26.375 173.830 ;
        RECT 25.335 173.220 26.375 173.390 ;
        RECT 26.590 173.360 26.760 173.690 ;
        RECT 27.100 172.820 27.390 174.230 ;
        RECT 24.440 172.700 27.390 172.820 ;
        RECT 24.440 172.650 27.270 172.700 ;
        RECT 14.430 172.250 17.260 172.300 ;
        RECT 14.310 172.130 17.260 172.250 ;
        RECT 14.310 170.720 14.600 172.130 ;
        RECT 14.940 171.260 15.110 171.590 ;
        RECT 15.325 171.560 16.365 171.730 ;
        RECT 15.325 171.120 16.365 171.290 ;
        RECT 16.580 171.260 16.750 171.590 ;
        RECT 17.090 170.720 17.260 172.130 ;
        RECT 14.310 170.600 17.260 170.720 ;
        RECT 14.430 170.550 17.260 170.600 ;
        RECT 17.820 172.220 20.560 172.290 ;
        RECT 21.140 172.220 23.880 172.290 ;
        RECT 17.820 172.120 20.690 172.220 ;
        RECT 17.820 170.710 17.990 172.120 ;
        RECT 18.330 171.250 18.500 171.580 ;
        RECT 18.670 171.550 19.710 171.720 ;
        RECT 18.670 171.110 19.710 171.280 ;
        RECT 19.880 171.250 20.050 171.580 ;
        RECT 20.390 170.710 20.690 172.120 ;
        RECT 17.820 170.570 20.690 170.710 ;
        RECT 21.010 172.120 23.880 172.220 ;
        RECT 21.010 170.710 21.310 172.120 ;
        RECT 21.650 171.250 21.820 171.580 ;
        RECT 21.990 171.550 23.030 171.720 ;
        RECT 21.990 171.110 23.030 171.280 ;
        RECT 23.200 171.250 23.370 171.580 ;
        RECT 23.710 170.710 23.880 172.120 ;
        RECT 21.010 170.570 23.880 170.710 ;
        RECT 17.820 170.540 20.560 170.570 ;
        RECT 21.140 170.540 23.880 170.570 ;
        RECT 24.440 172.250 27.270 172.300 ;
        RECT 24.440 172.130 27.390 172.250 ;
        RECT 24.440 170.720 24.610 172.130 ;
        RECT 24.950 171.260 25.120 171.590 ;
        RECT 25.335 171.560 26.375 171.730 ;
        RECT 25.335 171.120 26.375 171.290 ;
        RECT 26.590 171.260 26.760 171.590 ;
        RECT 27.100 170.720 27.390 172.130 ;
        RECT 24.440 170.600 27.390 170.720 ;
        RECT 24.440 170.550 27.270 170.600 ;
        RECT 14.430 170.150 17.260 170.200 ;
        RECT 14.310 170.030 17.260 170.150 ;
        RECT 14.310 168.620 14.600 170.030 ;
        RECT 14.940 169.160 15.110 169.490 ;
        RECT 15.325 169.460 16.365 169.630 ;
        RECT 15.325 169.020 16.365 169.190 ;
        RECT 16.580 169.160 16.750 169.490 ;
        RECT 17.090 168.620 17.260 170.030 ;
        RECT 14.310 168.500 17.260 168.620 ;
        RECT 14.430 168.450 17.260 168.500 ;
        RECT 17.820 170.120 20.560 170.190 ;
        RECT 21.140 170.120 23.880 170.190 ;
        RECT 17.820 170.020 20.690 170.120 ;
        RECT 17.820 168.610 17.990 170.020 ;
        RECT 18.330 169.150 18.500 169.480 ;
        RECT 18.670 169.450 19.710 169.620 ;
        RECT 18.670 169.010 19.710 169.180 ;
        RECT 19.880 169.150 20.050 169.480 ;
        RECT 20.390 168.610 20.690 170.020 ;
        RECT 17.820 168.470 20.690 168.610 ;
        RECT 21.010 170.020 23.880 170.120 ;
        RECT 21.010 168.610 21.310 170.020 ;
        RECT 21.650 169.150 21.820 169.480 ;
        RECT 21.990 169.450 23.030 169.620 ;
        RECT 21.990 169.010 23.030 169.180 ;
        RECT 23.200 169.150 23.370 169.480 ;
        RECT 23.710 168.610 23.880 170.020 ;
        RECT 21.010 168.470 23.880 168.610 ;
        RECT 17.820 168.440 20.560 168.470 ;
        RECT 21.140 168.440 23.880 168.470 ;
        RECT 24.440 170.150 27.270 170.200 ;
        RECT 24.440 170.030 27.390 170.150 ;
        RECT 24.440 168.620 24.610 170.030 ;
        RECT 24.950 169.160 25.120 169.490 ;
        RECT 25.335 169.460 26.375 169.630 ;
        RECT 25.335 169.020 26.375 169.190 ;
        RECT 26.590 169.160 26.760 169.490 ;
        RECT 27.100 168.620 27.390 170.030 ;
        RECT 24.440 168.500 27.390 168.620 ;
        RECT 24.440 168.450 27.270 168.500 ;
        RECT 14.430 168.050 17.260 168.100 ;
        RECT 14.310 167.930 17.260 168.050 ;
        RECT 14.310 166.520 14.600 167.930 ;
        RECT 14.940 167.060 15.110 167.390 ;
        RECT 15.325 167.360 16.365 167.530 ;
        RECT 15.325 166.920 16.365 167.090 ;
        RECT 16.580 167.060 16.750 167.390 ;
        RECT 17.090 166.520 17.260 167.930 ;
        RECT 14.310 166.400 17.260 166.520 ;
        RECT 14.430 166.350 17.260 166.400 ;
        RECT 17.820 168.020 20.560 168.090 ;
        RECT 21.140 168.020 23.880 168.090 ;
        RECT 17.820 167.920 20.690 168.020 ;
        RECT 17.820 166.510 17.990 167.920 ;
        RECT 18.330 167.050 18.500 167.380 ;
        RECT 18.670 167.350 19.710 167.520 ;
        RECT 18.670 166.910 19.710 167.080 ;
        RECT 19.880 167.050 20.050 167.380 ;
        RECT 20.390 166.510 20.690 167.920 ;
        RECT 17.820 166.370 20.690 166.510 ;
        RECT 21.010 167.920 23.880 168.020 ;
        RECT 21.010 166.510 21.310 167.920 ;
        RECT 21.650 167.050 21.820 167.380 ;
        RECT 21.990 167.350 23.030 167.520 ;
        RECT 21.990 166.910 23.030 167.080 ;
        RECT 23.200 167.050 23.370 167.380 ;
        RECT 23.710 166.510 23.880 167.920 ;
        RECT 21.010 166.370 23.880 166.510 ;
        RECT 17.820 166.340 20.560 166.370 ;
        RECT 21.140 166.340 23.880 166.370 ;
        RECT 24.440 168.050 27.270 168.100 ;
        RECT 24.440 167.930 27.390 168.050 ;
        RECT 24.440 166.520 24.610 167.930 ;
        RECT 24.950 167.060 25.120 167.390 ;
        RECT 25.335 167.360 26.375 167.530 ;
        RECT 25.335 166.920 26.375 167.090 ;
        RECT 26.590 167.060 26.760 167.390 ;
        RECT 27.100 166.520 27.390 167.930 ;
        RECT 24.440 166.400 27.390 166.520 ;
        RECT 24.440 166.350 27.270 166.400 ;
        RECT 14.430 165.950 17.260 166.000 ;
        RECT 14.310 165.830 17.260 165.950 ;
        RECT 14.310 164.420 14.600 165.830 ;
        RECT 14.940 164.960 15.110 165.290 ;
        RECT 15.325 165.260 16.365 165.430 ;
        RECT 15.325 164.820 16.365 164.990 ;
        RECT 16.580 164.960 16.750 165.290 ;
        RECT 17.090 164.420 17.260 165.830 ;
        RECT 14.310 164.300 17.260 164.420 ;
        RECT 14.430 164.250 17.260 164.300 ;
        RECT 17.820 165.920 20.560 165.990 ;
        RECT 21.140 165.920 23.880 165.990 ;
        RECT 17.820 165.820 20.690 165.920 ;
        RECT 17.820 164.410 17.990 165.820 ;
        RECT 18.330 164.950 18.500 165.280 ;
        RECT 18.670 165.250 19.710 165.420 ;
        RECT 18.670 164.810 19.710 164.980 ;
        RECT 19.880 164.950 20.050 165.280 ;
        RECT 20.390 164.410 20.690 165.820 ;
        RECT 17.820 164.270 20.690 164.410 ;
        RECT 21.010 165.820 23.880 165.920 ;
        RECT 21.010 164.410 21.310 165.820 ;
        RECT 21.650 164.950 21.820 165.280 ;
        RECT 21.990 165.250 23.030 165.420 ;
        RECT 21.990 164.810 23.030 164.980 ;
        RECT 23.200 164.950 23.370 165.280 ;
        RECT 23.710 164.410 23.880 165.820 ;
        RECT 21.010 164.270 23.880 164.410 ;
        RECT 17.820 164.240 20.560 164.270 ;
        RECT 21.140 164.240 23.880 164.270 ;
        RECT 24.440 165.950 27.270 166.000 ;
        RECT 24.440 165.830 27.390 165.950 ;
        RECT 24.440 164.420 24.610 165.830 ;
        RECT 24.950 164.960 25.120 165.290 ;
        RECT 25.335 165.260 26.375 165.430 ;
        RECT 25.335 164.820 26.375 164.990 ;
        RECT 26.590 164.960 26.760 165.290 ;
        RECT 27.100 164.420 27.390 165.830 ;
        RECT 24.440 164.300 27.390 164.420 ;
        RECT 24.440 164.250 27.270 164.300 ;
        RECT 14.430 163.850 17.260 163.900 ;
        RECT 14.310 163.730 17.260 163.850 ;
        RECT 14.310 162.320 14.600 163.730 ;
        RECT 14.940 162.860 15.110 163.190 ;
        RECT 15.325 163.160 16.365 163.330 ;
        RECT 15.325 162.720 16.365 162.890 ;
        RECT 16.580 162.860 16.750 163.190 ;
        RECT 17.090 162.320 17.260 163.730 ;
        RECT 14.310 162.200 17.260 162.320 ;
        RECT 14.430 162.150 17.260 162.200 ;
        RECT 17.820 163.820 20.560 163.890 ;
        RECT 21.140 163.820 23.880 163.890 ;
        RECT 17.820 163.720 20.690 163.820 ;
        RECT 17.820 162.310 17.990 163.720 ;
        RECT 18.330 162.850 18.500 163.180 ;
        RECT 18.670 163.150 19.710 163.320 ;
        RECT 18.670 162.710 19.710 162.880 ;
        RECT 19.880 162.850 20.050 163.180 ;
        RECT 20.390 162.310 20.690 163.720 ;
        RECT 17.820 162.170 20.690 162.310 ;
        RECT 21.010 163.720 23.880 163.820 ;
        RECT 21.010 162.310 21.310 163.720 ;
        RECT 21.650 162.850 21.820 163.180 ;
        RECT 21.990 163.150 23.030 163.320 ;
        RECT 21.990 162.710 23.030 162.880 ;
        RECT 23.200 162.850 23.370 163.180 ;
        RECT 23.710 162.310 23.880 163.720 ;
        RECT 21.010 162.170 23.880 162.310 ;
        RECT 17.820 162.140 20.560 162.170 ;
        RECT 21.140 162.140 23.880 162.170 ;
        RECT 24.440 163.850 27.270 163.900 ;
        RECT 24.440 163.730 27.390 163.850 ;
        RECT 24.440 162.320 24.610 163.730 ;
        RECT 24.950 162.860 25.120 163.190 ;
        RECT 25.335 163.160 26.375 163.330 ;
        RECT 25.335 162.720 26.375 162.890 ;
        RECT 26.590 162.860 26.760 163.190 ;
        RECT 27.100 162.320 27.390 163.730 ;
        RECT 24.440 162.200 27.390 162.320 ;
        RECT 24.440 162.150 27.270 162.200 ;
        RECT 14.430 161.750 17.260 161.800 ;
        RECT 14.310 161.630 17.260 161.750 ;
        RECT 14.310 160.220 14.600 161.630 ;
        RECT 14.940 160.760 15.110 161.090 ;
        RECT 15.325 161.060 16.365 161.230 ;
        RECT 15.325 160.620 16.365 160.790 ;
        RECT 16.580 160.760 16.750 161.090 ;
        RECT 17.090 160.220 17.260 161.630 ;
        RECT 14.310 160.100 17.260 160.220 ;
        RECT 14.430 160.050 17.260 160.100 ;
        RECT 17.820 161.720 20.560 161.790 ;
        RECT 21.140 161.720 23.880 161.790 ;
        RECT 17.820 161.620 20.690 161.720 ;
        RECT 17.820 160.210 17.990 161.620 ;
        RECT 18.330 160.750 18.500 161.080 ;
        RECT 18.670 161.050 19.710 161.220 ;
        RECT 18.670 160.610 19.710 160.780 ;
        RECT 19.880 160.750 20.050 161.080 ;
        RECT 20.390 160.210 20.690 161.620 ;
        RECT 17.820 160.070 20.690 160.210 ;
        RECT 21.010 161.620 23.880 161.720 ;
        RECT 21.010 160.210 21.310 161.620 ;
        RECT 21.650 160.750 21.820 161.080 ;
        RECT 21.990 161.050 23.030 161.220 ;
        RECT 21.990 160.610 23.030 160.780 ;
        RECT 23.200 160.750 23.370 161.080 ;
        RECT 23.710 160.210 23.880 161.620 ;
        RECT 21.010 160.070 23.880 160.210 ;
        RECT 17.820 160.040 20.560 160.070 ;
        RECT 21.140 160.040 23.880 160.070 ;
        RECT 24.440 161.750 27.270 161.800 ;
        RECT 24.440 161.630 27.390 161.750 ;
        RECT 24.440 160.220 24.610 161.630 ;
        RECT 24.950 160.760 25.120 161.090 ;
        RECT 25.335 161.060 26.375 161.230 ;
        RECT 25.335 160.620 26.375 160.790 ;
        RECT 26.590 160.760 26.760 161.090 ;
        RECT 27.100 160.220 27.390 161.630 ;
        RECT 24.440 160.100 27.390 160.220 ;
        RECT 24.440 160.050 27.270 160.100 ;
        RECT 14.430 159.650 17.260 159.700 ;
        RECT 14.310 159.530 17.260 159.650 ;
        RECT 14.310 158.120 14.600 159.530 ;
        RECT 14.940 158.660 15.110 158.990 ;
        RECT 15.325 158.960 16.365 159.130 ;
        RECT 15.325 158.520 16.365 158.690 ;
        RECT 16.580 158.660 16.750 158.990 ;
        RECT 17.090 158.120 17.260 159.530 ;
        RECT 14.310 158.000 17.260 158.120 ;
        RECT 14.430 157.950 17.260 158.000 ;
        RECT 17.820 159.620 20.560 159.690 ;
        RECT 21.140 159.620 23.880 159.690 ;
        RECT 17.820 159.520 20.690 159.620 ;
        RECT 17.820 158.110 17.990 159.520 ;
        RECT 18.330 158.650 18.500 158.980 ;
        RECT 18.670 158.950 19.710 159.120 ;
        RECT 18.670 158.510 19.710 158.680 ;
        RECT 19.880 158.650 20.050 158.980 ;
        RECT 20.390 158.110 20.690 159.520 ;
        RECT 17.820 157.970 20.690 158.110 ;
        RECT 21.010 159.520 23.880 159.620 ;
        RECT 21.010 158.110 21.310 159.520 ;
        RECT 21.650 158.650 21.820 158.980 ;
        RECT 21.990 158.950 23.030 159.120 ;
        RECT 21.990 158.510 23.030 158.680 ;
        RECT 23.200 158.650 23.370 158.980 ;
        RECT 23.710 158.110 23.880 159.520 ;
        RECT 21.010 157.970 23.880 158.110 ;
        RECT 17.820 157.940 20.560 157.970 ;
        RECT 21.140 157.940 23.880 157.970 ;
        RECT 24.440 159.650 27.270 159.700 ;
        RECT 24.440 159.530 27.390 159.650 ;
        RECT 24.440 158.120 24.610 159.530 ;
        RECT 24.950 158.660 25.120 158.990 ;
        RECT 25.335 158.960 26.375 159.130 ;
        RECT 25.335 158.520 26.375 158.690 ;
        RECT 26.590 158.660 26.760 158.990 ;
        RECT 27.100 158.120 27.390 159.530 ;
        RECT 24.440 158.000 27.390 158.120 ;
        RECT 24.440 157.950 27.270 158.000 ;
        RECT 14.430 157.550 17.260 157.600 ;
        RECT 14.310 157.430 17.260 157.550 ;
        RECT 14.310 156.020 14.600 157.430 ;
        RECT 14.940 156.560 15.110 156.890 ;
        RECT 15.325 156.860 16.365 157.030 ;
        RECT 15.325 156.420 16.365 156.590 ;
        RECT 16.580 156.560 16.750 156.890 ;
        RECT 17.090 156.020 17.260 157.430 ;
        RECT 14.310 155.900 17.260 156.020 ;
        RECT 14.430 155.850 17.260 155.900 ;
        RECT 17.820 157.520 20.560 157.590 ;
        RECT 21.140 157.520 23.880 157.590 ;
        RECT 17.820 157.420 20.690 157.520 ;
        RECT 17.820 156.010 17.990 157.420 ;
        RECT 18.330 156.550 18.500 156.880 ;
        RECT 18.670 156.850 19.710 157.020 ;
        RECT 18.670 156.410 19.710 156.580 ;
        RECT 19.880 156.550 20.050 156.880 ;
        RECT 20.390 156.010 20.690 157.420 ;
        RECT 17.820 155.870 20.690 156.010 ;
        RECT 21.010 157.420 23.880 157.520 ;
        RECT 21.010 156.010 21.310 157.420 ;
        RECT 21.650 156.550 21.820 156.880 ;
        RECT 21.990 156.850 23.030 157.020 ;
        RECT 21.990 156.410 23.030 156.580 ;
        RECT 23.200 156.550 23.370 156.880 ;
        RECT 23.710 156.010 23.880 157.420 ;
        RECT 21.010 155.870 23.880 156.010 ;
        RECT 17.820 155.840 20.560 155.870 ;
        RECT 21.140 155.840 23.880 155.870 ;
        RECT 24.440 157.550 27.270 157.600 ;
        RECT 24.440 157.430 27.390 157.550 ;
        RECT 24.440 156.020 24.610 157.430 ;
        RECT 24.950 156.560 25.120 156.890 ;
        RECT 25.335 156.860 26.375 157.030 ;
        RECT 25.335 156.420 26.375 156.590 ;
        RECT 26.590 156.560 26.760 156.890 ;
        RECT 27.100 156.020 27.390 157.430 ;
        RECT 24.440 155.900 27.390 156.020 ;
        RECT 24.440 155.850 27.270 155.900 ;
        RECT 14.430 155.450 17.260 155.500 ;
        RECT 14.310 155.330 17.260 155.450 ;
        RECT 14.310 153.920 14.600 155.330 ;
        RECT 14.940 154.460 15.110 154.790 ;
        RECT 15.325 154.760 16.365 154.930 ;
        RECT 15.325 154.320 16.365 154.490 ;
        RECT 16.580 154.460 16.750 154.790 ;
        RECT 17.090 153.920 17.260 155.330 ;
        RECT 14.310 153.800 17.260 153.920 ;
        RECT 14.430 153.750 17.260 153.800 ;
        RECT 17.820 155.420 20.560 155.490 ;
        RECT 21.140 155.420 23.880 155.490 ;
        RECT 17.820 155.320 20.690 155.420 ;
        RECT 17.820 153.910 17.990 155.320 ;
        RECT 18.330 154.450 18.500 154.780 ;
        RECT 18.670 154.750 19.710 154.920 ;
        RECT 18.670 154.310 19.710 154.480 ;
        RECT 19.880 154.450 20.050 154.780 ;
        RECT 20.390 153.910 20.690 155.320 ;
        RECT 17.820 153.770 20.690 153.910 ;
        RECT 21.010 155.320 23.880 155.420 ;
        RECT 21.010 153.910 21.310 155.320 ;
        RECT 21.650 154.450 21.820 154.780 ;
        RECT 21.990 154.750 23.030 154.920 ;
        RECT 21.990 154.310 23.030 154.480 ;
        RECT 23.200 154.450 23.370 154.780 ;
        RECT 23.710 153.910 23.880 155.320 ;
        RECT 21.010 153.770 23.880 153.910 ;
        RECT 17.820 153.740 20.560 153.770 ;
        RECT 21.140 153.740 23.880 153.770 ;
        RECT 24.440 155.450 27.270 155.500 ;
        RECT 24.440 155.330 27.390 155.450 ;
        RECT 24.440 153.920 24.610 155.330 ;
        RECT 24.950 154.460 25.120 154.790 ;
        RECT 25.335 154.760 26.375 154.930 ;
        RECT 25.335 154.320 26.375 154.490 ;
        RECT 26.590 154.460 26.760 154.790 ;
        RECT 27.100 153.920 27.390 155.330 ;
        RECT 24.440 153.800 27.390 153.920 ;
        RECT 24.440 153.750 27.270 153.800 ;
        RECT 14.430 153.350 17.260 153.400 ;
        RECT 14.310 153.230 17.260 153.350 ;
        RECT 14.310 151.820 14.600 153.230 ;
        RECT 14.940 152.360 15.110 152.690 ;
        RECT 15.325 152.660 16.365 152.830 ;
        RECT 15.325 152.220 16.365 152.390 ;
        RECT 16.580 152.360 16.750 152.690 ;
        RECT 17.090 151.820 17.260 153.230 ;
        RECT 14.310 151.700 17.260 151.820 ;
        RECT 14.430 151.650 17.260 151.700 ;
        RECT 17.820 153.320 20.560 153.390 ;
        RECT 21.140 153.320 23.880 153.390 ;
        RECT 17.820 153.220 20.690 153.320 ;
        RECT 17.820 151.810 17.990 153.220 ;
        RECT 18.330 152.350 18.500 152.680 ;
        RECT 18.670 152.650 19.710 152.820 ;
        RECT 18.670 152.210 19.710 152.380 ;
        RECT 19.880 152.350 20.050 152.680 ;
        RECT 20.390 151.810 20.690 153.220 ;
        RECT 17.820 151.670 20.690 151.810 ;
        RECT 21.010 153.220 23.880 153.320 ;
        RECT 21.010 151.810 21.310 153.220 ;
        RECT 21.650 152.350 21.820 152.680 ;
        RECT 21.990 152.650 23.030 152.820 ;
        RECT 21.990 152.210 23.030 152.380 ;
        RECT 23.200 152.350 23.370 152.680 ;
        RECT 23.710 151.810 23.880 153.220 ;
        RECT 21.010 151.670 23.880 151.810 ;
        RECT 17.820 151.640 20.560 151.670 ;
        RECT 21.140 151.640 23.880 151.670 ;
        RECT 24.440 153.350 27.270 153.400 ;
        RECT 24.440 153.230 27.390 153.350 ;
        RECT 24.440 151.820 24.610 153.230 ;
        RECT 24.950 152.360 25.120 152.690 ;
        RECT 25.335 152.660 26.375 152.830 ;
        RECT 25.335 152.220 26.375 152.390 ;
        RECT 26.590 152.360 26.760 152.690 ;
        RECT 27.100 151.820 27.390 153.230 ;
        RECT 24.440 151.700 27.390 151.820 ;
        RECT 24.440 151.650 27.270 151.700 ;
        RECT 14.430 151.250 17.260 151.300 ;
        RECT 14.310 151.130 17.260 151.250 ;
        RECT 14.310 149.720 14.600 151.130 ;
        RECT 14.940 150.260 15.110 150.590 ;
        RECT 15.325 150.560 16.365 150.730 ;
        RECT 15.325 150.120 16.365 150.290 ;
        RECT 16.580 150.260 16.750 150.590 ;
        RECT 17.090 149.720 17.260 151.130 ;
        RECT 14.310 149.600 17.260 149.720 ;
        RECT 14.430 149.550 17.260 149.600 ;
        RECT 17.820 151.220 20.560 151.290 ;
        RECT 21.140 151.220 23.880 151.290 ;
        RECT 17.820 151.120 20.690 151.220 ;
        RECT 17.820 149.710 17.990 151.120 ;
        RECT 18.330 150.250 18.500 150.580 ;
        RECT 18.670 150.550 19.710 150.720 ;
        RECT 18.670 150.110 19.710 150.280 ;
        RECT 19.880 150.250 20.050 150.580 ;
        RECT 20.390 149.710 20.690 151.120 ;
        RECT 17.820 149.570 20.690 149.710 ;
        RECT 21.010 151.120 23.880 151.220 ;
        RECT 21.010 149.710 21.310 151.120 ;
        RECT 21.650 150.250 21.820 150.580 ;
        RECT 21.990 150.550 23.030 150.720 ;
        RECT 21.990 150.110 23.030 150.280 ;
        RECT 23.200 150.250 23.370 150.580 ;
        RECT 23.710 149.710 23.880 151.120 ;
        RECT 21.010 149.570 23.880 149.710 ;
        RECT 17.820 149.540 20.560 149.570 ;
        RECT 21.140 149.540 23.880 149.570 ;
        RECT 24.440 151.250 27.270 151.300 ;
        RECT 24.440 151.130 27.390 151.250 ;
        RECT 24.440 149.720 24.610 151.130 ;
        RECT 24.950 150.260 25.120 150.590 ;
        RECT 25.335 150.560 26.375 150.730 ;
        RECT 25.335 150.120 26.375 150.290 ;
        RECT 26.590 150.260 26.760 150.590 ;
        RECT 27.100 149.720 27.390 151.130 ;
        RECT 24.440 149.600 27.390 149.720 ;
        RECT 24.440 149.550 27.270 149.600 ;
        RECT 14.430 149.150 17.260 149.200 ;
        RECT 14.310 149.030 17.260 149.150 ;
        RECT 14.310 147.620 14.600 149.030 ;
        RECT 14.940 148.160 15.110 148.490 ;
        RECT 15.325 148.460 16.365 148.630 ;
        RECT 15.325 148.020 16.365 148.190 ;
        RECT 16.580 148.160 16.750 148.490 ;
        RECT 17.090 147.620 17.260 149.030 ;
        RECT 14.310 147.500 17.260 147.620 ;
        RECT 14.430 147.450 17.260 147.500 ;
        RECT 17.820 149.120 20.560 149.190 ;
        RECT 21.140 149.120 23.880 149.190 ;
        RECT 17.820 149.020 20.690 149.120 ;
        RECT 17.820 147.610 17.990 149.020 ;
        RECT 18.330 148.150 18.500 148.480 ;
        RECT 18.670 148.450 19.710 148.620 ;
        RECT 18.670 148.010 19.710 148.180 ;
        RECT 19.880 148.150 20.050 148.480 ;
        RECT 20.390 147.610 20.690 149.020 ;
        RECT 17.820 147.470 20.690 147.610 ;
        RECT 21.010 149.020 23.880 149.120 ;
        RECT 21.010 147.610 21.310 149.020 ;
        RECT 21.650 148.150 21.820 148.480 ;
        RECT 21.990 148.450 23.030 148.620 ;
        RECT 21.990 148.010 23.030 148.180 ;
        RECT 23.200 148.150 23.370 148.480 ;
        RECT 23.710 147.610 23.880 149.020 ;
        RECT 21.010 147.470 23.880 147.610 ;
        RECT 17.820 147.440 20.560 147.470 ;
        RECT 21.140 147.440 23.880 147.470 ;
        RECT 24.440 149.150 27.270 149.200 ;
        RECT 24.440 149.030 27.390 149.150 ;
        RECT 24.440 147.620 24.610 149.030 ;
        RECT 24.950 148.160 25.120 148.490 ;
        RECT 25.335 148.460 26.375 148.630 ;
        RECT 25.335 148.020 26.375 148.190 ;
        RECT 26.590 148.160 26.760 148.490 ;
        RECT 27.100 147.620 27.390 149.030 ;
        RECT 24.440 147.500 27.390 147.620 ;
        RECT 24.440 147.450 27.270 147.500 ;
        RECT 14.430 147.050 17.260 147.100 ;
        RECT 14.310 146.930 17.260 147.050 ;
        RECT 14.310 145.520 14.600 146.930 ;
        RECT 14.940 146.060 15.110 146.390 ;
        RECT 15.325 146.360 16.365 146.530 ;
        RECT 15.325 145.920 16.365 146.090 ;
        RECT 16.580 146.060 16.750 146.390 ;
        RECT 17.090 145.520 17.260 146.930 ;
        RECT 14.310 145.400 17.260 145.520 ;
        RECT 14.430 145.350 17.260 145.400 ;
        RECT 17.820 147.020 20.560 147.090 ;
        RECT 21.140 147.020 23.880 147.090 ;
        RECT 17.820 146.920 20.690 147.020 ;
        RECT 17.820 145.510 17.990 146.920 ;
        RECT 18.330 146.050 18.500 146.380 ;
        RECT 18.670 146.350 19.710 146.520 ;
        RECT 18.670 145.910 19.710 146.080 ;
        RECT 19.880 146.050 20.050 146.380 ;
        RECT 20.390 145.510 20.690 146.920 ;
        RECT 17.820 145.370 20.690 145.510 ;
        RECT 21.010 146.920 23.880 147.020 ;
        RECT 21.010 145.510 21.310 146.920 ;
        RECT 21.650 146.050 21.820 146.380 ;
        RECT 21.990 146.350 23.030 146.520 ;
        RECT 21.990 145.910 23.030 146.080 ;
        RECT 23.200 146.050 23.370 146.380 ;
        RECT 23.710 145.510 23.880 146.920 ;
        RECT 21.010 145.370 23.880 145.510 ;
        RECT 17.820 145.340 20.560 145.370 ;
        RECT 21.140 145.340 23.880 145.370 ;
        RECT 24.440 147.050 27.270 147.100 ;
        RECT 24.440 146.930 27.390 147.050 ;
        RECT 24.440 145.520 24.610 146.930 ;
        RECT 24.950 146.060 25.120 146.390 ;
        RECT 25.335 146.360 26.375 146.530 ;
        RECT 25.335 145.920 26.375 146.090 ;
        RECT 26.590 146.060 26.760 146.390 ;
        RECT 27.100 145.520 27.390 146.930 ;
        RECT 24.440 145.400 27.390 145.520 ;
        RECT 24.440 145.350 27.270 145.400 ;
        RECT 14.430 144.950 17.260 145.000 ;
        RECT 14.310 144.830 17.260 144.950 ;
        RECT 14.310 143.420 14.600 144.830 ;
        RECT 14.940 143.960 15.110 144.290 ;
        RECT 15.325 144.260 16.365 144.430 ;
        RECT 15.325 143.820 16.365 143.990 ;
        RECT 16.580 143.960 16.750 144.290 ;
        RECT 17.090 143.420 17.260 144.830 ;
        RECT 14.310 143.300 17.260 143.420 ;
        RECT 14.430 143.250 17.260 143.300 ;
        RECT 17.820 144.920 20.560 144.990 ;
        RECT 21.140 144.920 23.880 144.990 ;
        RECT 17.820 144.820 20.690 144.920 ;
        RECT 17.820 143.410 17.990 144.820 ;
        RECT 18.330 143.950 18.500 144.280 ;
        RECT 18.670 144.250 19.710 144.420 ;
        RECT 18.670 143.810 19.710 143.980 ;
        RECT 19.880 143.950 20.050 144.280 ;
        RECT 20.390 143.410 20.690 144.820 ;
        RECT 17.820 143.270 20.690 143.410 ;
        RECT 21.010 144.820 23.880 144.920 ;
        RECT 21.010 143.410 21.310 144.820 ;
        RECT 21.650 143.950 21.820 144.280 ;
        RECT 21.990 144.250 23.030 144.420 ;
        RECT 21.990 143.810 23.030 143.980 ;
        RECT 23.200 143.950 23.370 144.280 ;
        RECT 23.710 143.410 23.880 144.820 ;
        RECT 21.010 143.270 23.880 143.410 ;
        RECT 17.820 143.240 20.560 143.270 ;
        RECT 21.140 143.240 23.880 143.270 ;
        RECT 24.440 144.950 27.270 145.000 ;
        RECT 24.440 144.830 27.390 144.950 ;
        RECT 24.440 143.420 24.610 144.830 ;
        RECT 24.950 143.960 25.120 144.290 ;
        RECT 25.335 144.260 26.375 144.430 ;
        RECT 25.335 143.820 26.375 143.990 ;
        RECT 26.590 143.960 26.760 144.290 ;
        RECT 27.100 143.420 27.390 144.830 ;
        RECT 24.440 143.300 27.390 143.420 ;
        RECT 24.440 143.250 27.270 143.300 ;
        RECT 14.430 142.850 17.260 142.900 ;
        RECT 14.310 142.730 17.260 142.850 ;
        RECT 14.310 141.320 14.600 142.730 ;
        RECT 14.940 141.860 15.110 142.190 ;
        RECT 15.325 142.160 16.365 142.330 ;
        RECT 15.325 141.720 16.365 141.890 ;
        RECT 16.580 141.860 16.750 142.190 ;
        RECT 17.090 141.320 17.260 142.730 ;
        RECT 14.310 141.200 17.260 141.320 ;
        RECT 14.430 141.150 17.260 141.200 ;
        RECT 17.820 142.820 20.560 142.890 ;
        RECT 21.140 142.820 23.880 142.890 ;
        RECT 17.820 142.720 20.690 142.820 ;
        RECT 17.820 141.310 17.990 142.720 ;
        RECT 18.330 141.850 18.500 142.180 ;
        RECT 18.670 142.150 19.710 142.320 ;
        RECT 18.670 141.710 19.710 141.880 ;
        RECT 19.880 141.850 20.050 142.180 ;
        RECT 20.390 141.310 20.690 142.720 ;
        RECT 17.820 141.170 20.690 141.310 ;
        RECT 21.010 142.720 23.880 142.820 ;
        RECT 21.010 141.310 21.310 142.720 ;
        RECT 21.650 141.850 21.820 142.180 ;
        RECT 21.990 142.150 23.030 142.320 ;
        RECT 21.990 141.710 23.030 141.880 ;
        RECT 23.200 141.850 23.370 142.180 ;
        RECT 23.710 141.310 23.880 142.720 ;
        RECT 21.010 141.170 23.880 141.310 ;
        RECT 17.820 141.140 20.560 141.170 ;
        RECT 21.140 141.140 23.880 141.170 ;
        RECT 24.440 142.850 27.270 142.900 ;
        RECT 24.440 142.730 27.390 142.850 ;
        RECT 24.440 141.320 24.610 142.730 ;
        RECT 24.950 141.860 25.120 142.190 ;
        RECT 25.335 142.160 26.375 142.330 ;
        RECT 25.335 141.720 26.375 141.890 ;
        RECT 26.590 141.860 26.760 142.190 ;
        RECT 27.100 141.320 27.390 142.730 ;
        RECT 24.440 141.200 27.390 141.320 ;
        RECT 24.440 141.150 27.270 141.200 ;
        RECT 14.430 140.750 17.260 140.800 ;
        RECT 14.310 140.630 17.260 140.750 ;
        RECT 14.310 139.220 14.600 140.630 ;
        RECT 14.940 139.760 15.110 140.090 ;
        RECT 15.325 140.060 16.365 140.230 ;
        RECT 15.325 139.620 16.365 139.790 ;
        RECT 16.580 139.760 16.750 140.090 ;
        RECT 17.090 139.220 17.260 140.630 ;
        RECT 14.310 139.100 17.260 139.220 ;
        RECT 14.430 139.050 17.260 139.100 ;
        RECT 17.820 140.720 20.560 140.790 ;
        RECT 21.140 140.720 23.880 140.790 ;
        RECT 17.820 140.620 20.690 140.720 ;
        RECT 17.820 139.210 17.990 140.620 ;
        RECT 18.330 139.750 18.500 140.080 ;
        RECT 18.670 140.050 19.710 140.220 ;
        RECT 18.670 139.610 19.710 139.780 ;
        RECT 19.880 139.750 20.050 140.080 ;
        RECT 20.390 139.210 20.690 140.620 ;
        RECT 17.820 139.070 20.690 139.210 ;
        RECT 21.010 140.620 23.880 140.720 ;
        RECT 21.010 139.210 21.310 140.620 ;
        RECT 21.650 139.750 21.820 140.080 ;
        RECT 21.990 140.050 23.030 140.220 ;
        RECT 21.990 139.610 23.030 139.780 ;
        RECT 23.200 139.750 23.370 140.080 ;
        RECT 23.710 139.210 23.880 140.620 ;
        RECT 21.010 139.070 23.880 139.210 ;
        RECT 17.820 139.040 20.560 139.070 ;
        RECT 21.140 139.040 23.880 139.070 ;
        RECT 24.440 140.750 27.270 140.800 ;
        RECT 24.440 140.630 27.390 140.750 ;
        RECT 24.440 139.220 24.610 140.630 ;
        RECT 24.950 139.760 25.120 140.090 ;
        RECT 25.335 140.060 26.375 140.230 ;
        RECT 25.335 139.620 26.375 139.790 ;
        RECT 26.590 139.760 26.760 140.090 ;
        RECT 27.100 139.220 27.390 140.630 ;
        RECT 24.440 139.100 27.390 139.220 ;
        RECT 24.440 139.050 27.270 139.100 ;
        RECT 14.430 138.650 17.260 138.700 ;
        RECT 14.310 138.530 17.260 138.650 ;
        RECT 14.310 137.120 14.600 138.530 ;
        RECT 14.940 137.660 15.110 137.990 ;
        RECT 15.325 137.960 16.365 138.130 ;
        RECT 15.325 137.520 16.365 137.690 ;
        RECT 16.580 137.660 16.750 137.990 ;
        RECT 17.090 137.120 17.260 138.530 ;
        RECT 14.310 137.000 17.260 137.120 ;
        RECT 14.430 136.950 17.260 137.000 ;
        RECT 17.820 138.620 20.560 138.690 ;
        RECT 21.140 138.620 23.880 138.690 ;
        RECT 17.820 138.520 20.690 138.620 ;
        RECT 17.820 137.110 17.990 138.520 ;
        RECT 18.330 137.650 18.500 137.980 ;
        RECT 18.670 137.950 19.710 138.120 ;
        RECT 18.670 137.510 19.710 137.680 ;
        RECT 19.880 137.650 20.050 137.980 ;
        RECT 20.390 137.110 20.690 138.520 ;
        RECT 17.820 136.970 20.690 137.110 ;
        RECT 21.010 138.520 23.880 138.620 ;
        RECT 21.010 137.110 21.310 138.520 ;
        RECT 21.650 137.650 21.820 137.980 ;
        RECT 21.990 137.950 23.030 138.120 ;
        RECT 21.990 137.510 23.030 137.680 ;
        RECT 23.200 137.650 23.370 137.980 ;
        RECT 23.710 137.110 23.880 138.520 ;
        RECT 21.010 136.970 23.880 137.110 ;
        RECT 17.820 136.940 20.560 136.970 ;
        RECT 21.140 136.940 23.880 136.970 ;
        RECT 24.440 138.650 27.270 138.700 ;
        RECT 24.440 138.530 27.390 138.650 ;
        RECT 24.440 137.120 24.610 138.530 ;
        RECT 24.950 137.660 25.120 137.990 ;
        RECT 25.335 137.960 26.375 138.130 ;
        RECT 25.335 137.520 26.375 137.690 ;
        RECT 26.590 137.660 26.760 137.990 ;
        RECT 27.100 137.120 27.390 138.530 ;
        RECT 24.440 137.000 27.390 137.120 ;
        RECT 24.440 136.950 27.270 137.000 ;
        RECT 14.430 136.550 17.260 136.600 ;
        RECT 14.310 136.430 17.260 136.550 ;
        RECT 14.310 135.020 14.600 136.430 ;
        RECT 14.940 135.560 15.110 135.890 ;
        RECT 15.325 135.860 16.365 136.030 ;
        RECT 15.325 135.420 16.365 135.590 ;
        RECT 16.580 135.560 16.750 135.890 ;
        RECT 17.090 135.020 17.260 136.430 ;
        RECT 14.310 134.900 17.260 135.020 ;
        RECT 14.430 134.850 17.260 134.900 ;
        RECT 17.820 136.520 20.560 136.590 ;
        RECT 21.140 136.520 23.880 136.590 ;
        RECT 17.820 136.420 20.690 136.520 ;
        RECT 17.820 135.010 17.990 136.420 ;
        RECT 18.330 135.550 18.500 135.880 ;
        RECT 18.670 135.850 19.710 136.020 ;
        RECT 18.670 135.410 19.710 135.580 ;
        RECT 19.880 135.550 20.050 135.880 ;
        RECT 20.390 135.010 20.690 136.420 ;
        RECT 17.820 134.870 20.690 135.010 ;
        RECT 21.010 136.420 23.880 136.520 ;
        RECT 21.010 135.010 21.310 136.420 ;
        RECT 21.650 135.550 21.820 135.880 ;
        RECT 21.990 135.850 23.030 136.020 ;
        RECT 21.990 135.410 23.030 135.580 ;
        RECT 23.200 135.550 23.370 135.880 ;
        RECT 23.710 135.010 23.880 136.420 ;
        RECT 21.010 134.870 23.880 135.010 ;
        RECT 17.820 134.840 20.560 134.870 ;
        RECT 21.140 134.840 23.880 134.870 ;
        RECT 24.440 136.550 27.270 136.600 ;
        RECT 24.440 136.430 27.390 136.550 ;
        RECT 24.440 135.020 24.610 136.430 ;
        RECT 24.950 135.560 25.120 135.890 ;
        RECT 25.335 135.860 26.375 136.030 ;
        RECT 25.335 135.420 26.375 135.590 ;
        RECT 26.590 135.560 26.760 135.890 ;
        RECT 27.100 135.020 27.390 136.430 ;
        RECT 24.440 134.900 27.390 135.020 ;
        RECT 24.440 134.850 27.270 134.900 ;
        RECT 14.430 134.450 17.260 134.500 ;
        RECT 14.310 134.330 17.260 134.450 ;
        RECT 14.310 132.920 14.600 134.330 ;
        RECT 14.940 133.460 15.110 133.790 ;
        RECT 15.325 133.760 16.365 133.930 ;
        RECT 15.325 133.320 16.365 133.490 ;
        RECT 16.580 133.460 16.750 133.790 ;
        RECT 17.090 132.920 17.260 134.330 ;
        RECT 14.310 132.800 17.260 132.920 ;
        RECT 14.430 132.750 17.260 132.800 ;
        RECT 17.820 134.420 20.560 134.490 ;
        RECT 21.140 134.420 23.880 134.490 ;
        RECT 17.820 134.320 20.690 134.420 ;
        RECT 17.820 132.910 17.990 134.320 ;
        RECT 18.330 133.450 18.500 133.780 ;
        RECT 18.670 133.750 19.710 133.920 ;
        RECT 18.670 133.310 19.710 133.480 ;
        RECT 19.880 133.450 20.050 133.780 ;
        RECT 20.390 132.910 20.690 134.320 ;
        RECT 17.820 132.770 20.690 132.910 ;
        RECT 21.010 134.320 23.880 134.420 ;
        RECT 21.010 132.910 21.310 134.320 ;
        RECT 21.650 133.450 21.820 133.780 ;
        RECT 21.990 133.750 23.030 133.920 ;
        RECT 21.990 133.310 23.030 133.480 ;
        RECT 23.200 133.450 23.370 133.780 ;
        RECT 23.710 132.910 23.880 134.320 ;
        RECT 21.010 132.770 23.880 132.910 ;
        RECT 17.820 132.740 20.560 132.770 ;
        RECT 21.140 132.740 23.880 132.770 ;
        RECT 24.440 134.450 27.270 134.500 ;
        RECT 24.440 134.330 27.390 134.450 ;
        RECT 24.440 132.920 24.610 134.330 ;
        RECT 24.950 133.460 25.120 133.790 ;
        RECT 25.335 133.760 26.375 133.930 ;
        RECT 25.335 133.320 26.375 133.490 ;
        RECT 26.590 133.460 26.760 133.790 ;
        RECT 27.100 132.920 27.390 134.330 ;
        RECT 24.440 132.800 27.390 132.920 ;
        RECT 24.440 132.750 27.270 132.800 ;
        RECT 14.430 132.350 17.260 132.400 ;
        RECT 14.310 132.230 17.260 132.350 ;
        RECT 14.310 130.820 14.600 132.230 ;
        RECT 14.940 131.360 15.110 131.690 ;
        RECT 15.325 131.660 16.365 131.830 ;
        RECT 15.325 131.220 16.365 131.390 ;
        RECT 16.580 131.360 16.750 131.690 ;
        RECT 17.090 130.820 17.260 132.230 ;
        RECT 14.310 130.700 17.260 130.820 ;
        RECT 14.430 130.650 17.260 130.700 ;
        RECT 17.820 132.320 20.560 132.390 ;
        RECT 21.140 132.320 23.880 132.390 ;
        RECT 17.820 132.220 20.690 132.320 ;
        RECT 17.820 130.810 17.990 132.220 ;
        RECT 18.330 131.350 18.500 131.680 ;
        RECT 18.670 131.650 19.710 131.820 ;
        RECT 18.670 131.210 19.710 131.380 ;
        RECT 19.880 131.350 20.050 131.680 ;
        RECT 20.390 130.810 20.690 132.220 ;
        RECT 17.820 130.670 20.690 130.810 ;
        RECT 21.010 132.220 23.880 132.320 ;
        RECT 21.010 130.810 21.310 132.220 ;
        RECT 21.650 131.350 21.820 131.680 ;
        RECT 21.990 131.650 23.030 131.820 ;
        RECT 21.990 131.210 23.030 131.380 ;
        RECT 23.200 131.350 23.370 131.680 ;
        RECT 23.710 130.810 23.880 132.220 ;
        RECT 21.010 130.670 23.880 130.810 ;
        RECT 17.820 130.640 20.560 130.670 ;
        RECT 21.140 130.640 23.880 130.670 ;
        RECT 24.440 132.350 27.270 132.400 ;
        RECT 24.440 132.230 27.390 132.350 ;
        RECT 24.440 130.820 24.610 132.230 ;
        RECT 24.950 131.360 25.120 131.690 ;
        RECT 25.335 131.660 26.375 131.830 ;
        RECT 25.335 131.220 26.375 131.390 ;
        RECT 26.590 131.360 26.760 131.690 ;
        RECT 27.100 130.820 27.390 132.230 ;
        RECT 24.440 130.700 27.390 130.820 ;
        RECT 24.440 130.650 27.270 130.700 ;
        RECT 14.430 130.250 17.260 130.300 ;
        RECT 14.310 130.130 17.260 130.250 ;
        RECT 14.310 128.720 14.600 130.130 ;
        RECT 14.940 129.260 15.110 129.590 ;
        RECT 15.325 129.560 16.365 129.730 ;
        RECT 15.325 129.120 16.365 129.290 ;
        RECT 16.580 129.260 16.750 129.590 ;
        RECT 17.090 128.720 17.260 130.130 ;
        RECT 14.310 128.600 17.260 128.720 ;
        RECT 14.430 128.550 17.260 128.600 ;
        RECT 17.820 130.220 20.560 130.290 ;
        RECT 21.140 130.220 23.880 130.290 ;
        RECT 17.820 130.120 20.690 130.220 ;
        RECT 17.820 128.710 17.990 130.120 ;
        RECT 18.330 129.250 18.500 129.580 ;
        RECT 18.670 129.550 19.710 129.720 ;
        RECT 18.670 129.110 19.710 129.280 ;
        RECT 19.880 129.250 20.050 129.580 ;
        RECT 20.390 128.710 20.690 130.120 ;
        RECT 17.820 128.570 20.690 128.710 ;
        RECT 21.010 130.120 23.880 130.220 ;
        RECT 21.010 128.710 21.310 130.120 ;
        RECT 21.650 129.250 21.820 129.580 ;
        RECT 21.990 129.550 23.030 129.720 ;
        RECT 21.990 129.110 23.030 129.280 ;
        RECT 23.200 129.250 23.370 129.580 ;
        RECT 23.710 128.710 23.880 130.120 ;
        RECT 21.010 128.570 23.880 128.710 ;
        RECT 17.820 128.540 20.560 128.570 ;
        RECT 21.140 128.540 23.880 128.570 ;
        RECT 24.440 130.250 27.270 130.300 ;
        RECT 24.440 130.130 27.390 130.250 ;
        RECT 24.440 128.720 24.610 130.130 ;
        RECT 24.950 129.260 25.120 129.590 ;
        RECT 25.335 129.560 26.375 129.730 ;
        RECT 25.335 129.120 26.375 129.290 ;
        RECT 26.590 129.260 26.760 129.590 ;
        RECT 27.100 128.720 27.390 130.130 ;
        RECT 24.440 128.600 27.390 128.720 ;
        RECT 24.440 128.550 27.270 128.600 ;
        RECT 14.430 128.150 17.260 128.200 ;
        RECT 14.310 128.030 17.260 128.150 ;
        RECT 14.310 126.620 14.600 128.030 ;
        RECT 14.940 127.160 15.110 127.490 ;
        RECT 15.325 127.460 16.365 127.630 ;
        RECT 15.325 127.020 16.365 127.190 ;
        RECT 16.580 127.160 16.750 127.490 ;
        RECT 17.090 126.620 17.260 128.030 ;
        RECT 14.310 126.500 17.260 126.620 ;
        RECT 14.430 126.450 17.260 126.500 ;
        RECT 17.820 128.120 20.560 128.190 ;
        RECT 21.140 128.120 23.880 128.190 ;
        RECT 17.820 128.020 20.690 128.120 ;
        RECT 17.820 126.610 17.990 128.020 ;
        RECT 18.330 127.150 18.500 127.480 ;
        RECT 18.670 127.450 19.710 127.620 ;
        RECT 18.670 127.010 19.710 127.180 ;
        RECT 19.880 127.150 20.050 127.480 ;
        RECT 20.390 126.610 20.690 128.020 ;
        RECT 17.820 126.470 20.690 126.610 ;
        RECT 21.010 128.020 23.880 128.120 ;
        RECT 21.010 126.610 21.310 128.020 ;
        RECT 21.650 127.150 21.820 127.480 ;
        RECT 21.990 127.450 23.030 127.620 ;
        RECT 21.990 127.010 23.030 127.180 ;
        RECT 23.200 127.150 23.370 127.480 ;
        RECT 23.710 126.610 23.880 128.020 ;
        RECT 21.010 126.470 23.880 126.610 ;
        RECT 17.820 126.440 20.560 126.470 ;
        RECT 21.140 126.440 23.880 126.470 ;
        RECT 24.440 128.150 27.270 128.200 ;
        RECT 24.440 128.030 27.390 128.150 ;
        RECT 24.440 126.620 24.610 128.030 ;
        RECT 24.950 127.160 25.120 127.490 ;
        RECT 25.335 127.460 26.375 127.630 ;
        RECT 25.335 127.020 26.375 127.190 ;
        RECT 26.590 127.160 26.760 127.490 ;
        RECT 27.100 126.620 27.390 128.030 ;
        RECT 24.440 126.500 27.390 126.620 ;
        RECT 24.440 126.450 27.270 126.500 ;
        RECT 14.430 126.050 17.260 126.100 ;
        RECT 14.310 125.930 17.260 126.050 ;
        RECT 14.310 124.520 14.600 125.930 ;
        RECT 14.940 125.060 15.110 125.390 ;
        RECT 15.325 125.360 16.365 125.530 ;
        RECT 15.325 124.920 16.365 125.090 ;
        RECT 16.580 125.060 16.750 125.390 ;
        RECT 17.090 124.520 17.260 125.930 ;
        RECT 14.310 124.400 17.260 124.520 ;
        RECT 14.430 124.350 17.260 124.400 ;
        RECT 17.820 126.020 20.560 126.090 ;
        RECT 21.140 126.020 23.880 126.090 ;
        RECT 17.820 125.920 20.690 126.020 ;
        RECT 17.820 124.510 17.990 125.920 ;
        RECT 18.330 125.050 18.500 125.380 ;
        RECT 18.670 125.350 19.710 125.520 ;
        RECT 18.670 124.910 19.710 125.080 ;
        RECT 19.880 125.050 20.050 125.380 ;
        RECT 20.390 124.510 20.690 125.920 ;
        RECT 17.820 124.370 20.690 124.510 ;
        RECT 21.010 125.920 23.880 126.020 ;
        RECT 21.010 124.510 21.310 125.920 ;
        RECT 21.650 125.050 21.820 125.380 ;
        RECT 21.990 125.350 23.030 125.520 ;
        RECT 21.990 124.910 23.030 125.080 ;
        RECT 23.200 125.050 23.370 125.380 ;
        RECT 23.710 124.510 23.880 125.920 ;
        RECT 21.010 124.370 23.880 124.510 ;
        RECT 17.820 124.340 20.560 124.370 ;
        RECT 21.140 124.340 23.880 124.370 ;
        RECT 24.440 126.050 27.270 126.100 ;
        RECT 24.440 125.930 27.390 126.050 ;
        RECT 24.440 124.520 24.610 125.930 ;
        RECT 24.950 125.060 25.120 125.390 ;
        RECT 25.335 125.360 26.375 125.530 ;
        RECT 25.335 124.920 26.375 125.090 ;
        RECT 26.590 125.060 26.760 125.390 ;
        RECT 27.100 124.520 27.390 125.930 ;
        RECT 24.440 124.400 27.390 124.520 ;
        RECT 24.440 124.350 27.270 124.400 ;
        RECT 14.430 123.950 17.260 124.000 ;
        RECT 14.310 123.830 17.260 123.950 ;
        RECT 14.310 122.420 14.600 123.830 ;
        RECT 14.940 122.960 15.110 123.290 ;
        RECT 15.325 123.260 16.365 123.430 ;
        RECT 15.325 122.820 16.365 122.990 ;
        RECT 16.580 122.960 16.750 123.290 ;
        RECT 17.090 122.420 17.260 123.830 ;
        RECT 14.310 122.300 17.260 122.420 ;
        RECT 14.430 122.250 17.260 122.300 ;
        RECT 17.820 123.920 20.560 123.990 ;
        RECT 21.140 123.920 23.880 123.990 ;
        RECT 17.820 123.820 20.690 123.920 ;
        RECT 17.820 122.410 17.990 123.820 ;
        RECT 18.330 122.950 18.500 123.280 ;
        RECT 18.670 123.250 19.710 123.420 ;
        RECT 18.670 122.810 19.710 122.980 ;
        RECT 19.880 122.950 20.050 123.280 ;
        RECT 20.390 122.410 20.690 123.820 ;
        RECT 17.820 122.270 20.690 122.410 ;
        RECT 21.010 123.820 23.880 123.920 ;
        RECT 21.010 122.410 21.310 123.820 ;
        RECT 21.650 122.950 21.820 123.280 ;
        RECT 21.990 123.250 23.030 123.420 ;
        RECT 21.990 122.810 23.030 122.980 ;
        RECT 23.200 122.950 23.370 123.280 ;
        RECT 23.710 122.410 23.880 123.820 ;
        RECT 21.010 122.270 23.880 122.410 ;
        RECT 17.820 122.240 20.560 122.270 ;
        RECT 21.140 122.240 23.880 122.270 ;
        RECT 24.440 123.950 27.270 124.000 ;
        RECT 24.440 123.830 27.390 123.950 ;
        RECT 24.440 122.420 24.610 123.830 ;
        RECT 24.950 122.960 25.120 123.290 ;
        RECT 25.335 123.260 26.375 123.430 ;
        RECT 25.335 122.820 26.375 122.990 ;
        RECT 26.590 122.960 26.760 123.290 ;
        RECT 27.100 122.420 27.390 123.830 ;
        RECT 24.440 122.300 27.390 122.420 ;
        RECT 24.440 122.250 27.270 122.300 ;
        RECT 14.430 121.850 17.260 121.900 ;
        RECT 14.310 121.730 17.260 121.850 ;
        RECT 14.310 120.320 14.600 121.730 ;
        RECT 14.940 120.860 15.110 121.190 ;
        RECT 15.325 121.160 16.365 121.330 ;
        RECT 15.325 120.720 16.365 120.890 ;
        RECT 16.580 120.860 16.750 121.190 ;
        RECT 17.090 120.320 17.260 121.730 ;
        RECT 14.310 120.200 17.260 120.320 ;
        RECT 14.430 120.150 17.260 120.200 ;
        RECT 17.820 121.820 20.560 121.890 ;
        RECT 21.140 121.820 23.880 121.890 ;
        RECT 17.820 121.720 20.690 121.820 ;
        RECT 17.820 120.310 17.990 121.720 ;
        RECT 18.330 120.850 18.500 121.180 ;
        RECT 18.670 121.150 19.710 121.320 ;
        RECT 18.670 120.710 19.710 120.880 ;
        RECT 19.880 120.850 20.050 121.180 ;
        RECT 20.390 120.310 20.690 121.720 ;
        RECT 17.820 120.170 20.690 120.310 ;
        RECT 21.010 121.720 23.880 121.820 ;
        RECT 21.010 120.310 21.310 121.720 ;
        RECT 21.650 120.850 21.820 121.180 ;
        RECT 21.990 121.150 23.030 121.320 ;
        RECT 21.990 120.710 23.030 120.880 ;
        RECT 23.200 120.850 23.370 121.180 ;
        RECT 23.710 120.310 23.880 121.720 ;
        RECT 21.010 120.170 23.880 120.310 ;
        RECT 17.820 120.140 20.560 120.170 ;
        RECT 21.140 120.140 23.880 120.170 ;
        RECT 24.440 121.850 27.270 121.900 ;
        RECT 24.440 121.730 27.390 121.850 ;
        RECT 24.440 120.320 24.610 121.730 ;
        RECT 24.950 120.860 25.120 121.190 ;
        RECT 25.335 121.160 26.375 121.330 ;
        RECT 25.335 120.720 26.375 120.890 ;
        RECT 26.590 120.860 26.760 121.190 ;
        RECT 27.100 120.320 27.390 121.730 ;
        RECT 24.440 120.200 27.390 120.320 ;
        RECT 24.440 120.150 27.270 120.200 ;
        RECT 14.430 119.750 17.260 119.800 ;
        RECT 14.310 119.630 17.260 119.750 ;
        RECT 14.310 118.220 14.600 119.630 ;
        RECT 14.940 118.760 15.110 119.090 ;
        RECT 15.325 119.060 16.365 119.230 ;
        RECT 15.325 118.620 16.365 118.790 ;
        RECT 16.580 118.760 16.750 119.090 ;
        RECT 17.090 118.220 17.260 119.630 ;
        RECT 14.310 118.100 17.260 118.220 ;
        RECT 14.430 118.050 17.260 118.100 ;
        RECT 17.820 119.720 20.560 119.790 ;
        RECT 21.140 119.720 23.880 119.790 ;
        RECT 17.820 119.620 20.690 119.720 ;
        RECT 17.820 118.210 17.990 119.620 ;
        RECT 18.330 118.750 18.500 119.080 ;
        RECT 18.670 119.050 19.710 119.220 ;
        RECT 18.670 118.610 19.710 118.780 ;
        RECT 19.880 118.750 20.050 119.080 ;
        RECT 20.390 118.210 20.690 119.620 ;
        RECT 17.820 118.070 20.690 118.210 ;
        RECT 21.010 119.620 23.880 119.720 ;
        RECT 21.010 118.210 21.310 119.620 ;
        RECT 21.650 118.750 21.820 119.080 ;
        RECT 21.990 119.050 23.030 119.220 ;
        RECT 21.990 118.610 23.030 118.780 ;
        RECT 23.200 118.750 23.370 119.080 ;
        RECT 23.710 118.210 23.880 119.620 ;
        RECT 21.010 118.070 23.880 118.210 ;
        RECT 17.820 118.040 20.560 118.070 ;
        RECT 21.140 118.040 23.880 118.070 ;
        RECT 24.440 119.750 27.270 119.800 ;
        RECT 24.440 119.630 27.390 119.750 ;
        RECT 24.440 118.220 24.610 119.630 ;
        RECT 24.950 118.760 25.120 119.090 ;
        RECT 25.335 119.060 26.375 119.230 ;
        RECT 25.335 118.620 26.375 118.790 ;
        RECT 26.590 118.760 26.760 119.090 ;
        RECT 27.100 118.220 27.390 119.630 ;
        RECT 24.440 118.100 27.390 118.220 ;
        RECT 24.440 118.050 27.270 118.100 ;
        RECT 14.430 117.650 17.260 117.700 ;
        RECT 14.310 117.530 17.260 117.650 ;
        RECT 14.310 116.120 14.600 117.530 ;
        RECT 14.940 116.660 15.110 116.990 ;
        RECT 15.325 116.960 16.365 117.130 ;
        RECT 15.325 116.520 16.365 116.690 ;
        RECT 16.580 116.660 16.750 116.990 ;
        RECT 17.090 116.120 17.260 117.530 ;
        RECT 14.310 116.000 17.260 116.120 ;
        RECT 14.430 115.950 17.260 116.000 ;
        RECT 17.820 117.620 20.560 117.690 ;
        RECT 21.140 117.620 23.880 117.690 ;
        RECT 17.820 117.520 20.690 117.620 ;
        RECT 17.820 116.110 17.990 117.520 ;
        RECT 18.330 116.650 18.500 116.980 ;
        RECT 18.670 116.950 19.710 117.120 ;
        RECT 18.670 116.510 19.710 116.680 ;
        RECT 19.880 116.650 20.050 116.980 ;
        RECT 20.390 116.110 20.690 117.520 ;
        RECT 17.820 115.970 20.690 116.110 ;
        RECT 21.010 117.520 23.880 117.620 ;
        RECT 21.010 116.110 21.310 117.520 ;
        RECT 21.650 116.650 21.820 116.980 ;
        RECT 21.990 116.950 23.030 117.120 ;
        RECT 21.990 116.510 23.030 116.680 ;
        RECT 23.200 116.650 23.370 116.980 ;
        RECT 23.710 116.110 23.880 117.520 ;
        RECT 21.010 115.970 23.880 116.110 ;
        RECT 17.820 115.940 20.560 115.970 ;
        RECT 21.140 115.940 23.880 115.970 ;
        RECT 24.440 117.650 27.270 117.700 ;
        RECT 24.440 117.530 27.390 117.650 ;
        RECT 24.440 116.120 24.610 117.530 ;
        RECT 24.950 116.660 25.120 116.990 ;
        RECT 25.335 116.960 26.375 117.130 ;
        RECT 25.335 116.520 26.375 116.690 ;
        RECT 26.590 116.660 26.760 116.990 ;
        RECT 27.100 116.120 27.390 117.530 ;
        RECT 24.440 116.000 27.390 116.120 ;
        RECT 24.440 115.950 27.270 116.000 ;
        RECT 14.430 115.550 17.260 115.600 ;
        RECT 14.310 115.430 17.260 115.550 ;
        RECT 14.310 114.020 14.600 115.430 ;
        RECT 14.940 114.560 15.110 114.890 ;
        RECT 15.325 114.860 16.365 115.030 ;
        RECT 15.325 114.420 16.365 114.590 ;
        RECT 16.580 114.560 16.750 114.890 ;
        RECT 17.090 114.020 17.260 115.430 ;
        RECT 14.310 113.900 17.260 114.020 ;
        RECT 14.430 113.850 17.260 113.900 ;
        RECT 17.820 115.520 20.560 115.590 ;
        RECT 21.140 115.520 23.880 115.590 ;
        RECT 17.820 115.420 20.690 115.520 ;
        RECT 17.820 114.010 17.990 115.420 ;
        RECT 18.330 114.550 18.500 114.880 ;
        RECT 18.670 114.850 19.710 115.020 ;
        RECT 18.670 114.410 19.710 114.580 ;
        RECT 19.880 114.550 20.050 114.880 ;
        RECT 20.390 114.010 20.690 115.420 ;
        RECT 17.820 113.870 20.690 114.010 ;
        RECT 21.010 115.420 23.880 115.520 ;
        RECT 21.010 114.010 21.310 115.420 ;
        RECT 21.650 114.550 21.820 114.880 ;
        RECT 21.990 114.850 23.030 115.020 ;
        RECT 21.990 114.410 23.030 114.580 ;
        RECT 23.200 114.550 23.370 114.880 ;
        RECT 23.710 114.010 23.880 115.420 ;
        RECT 21.010 113.870 23.880 114.010 ;
        RECT 17.820 113.840 20.560 113.870 ;
        RECT 21.140 113.840 23.880 113.870 ;
        RECT 24.440 115.550 27.270 115.600 ;
        RECT 24.440 115.430 27.390 115.550 ;
        RECT 24.440 114.020 24.610 115.430 ;
        RECT 24.950 114.560 25.120 114.890 ;
        RECT 25.335 114.860 26.375 115.030 ;
        RECT 25.335 114.420 26.375 114.590 ;
        RECT 26.590 114.560 26.760 114.890 ;
        RECT 27.100 114.020 27.390 115.430 ;
        RECT 24.440 113.900 27.390 114.020 ;
        RECT 24.440 113.850 27.270 113.900 ;
        RECT 14.430 113.450 17.260 113.500 ;
        RECT 14.310 113.330 17.260 113.450 ;
        RECT 14.310 111.920 14.600 113.330 ;
        RECT 14.940 112.460 15.110 112.790 ;
        RECT 15.325 112.760 16.365 112.930 ;
        RECT 15.325 112.320 16.365 112.490 ;
        RECT 16.580 112.460 16.750 112.790 ;
        RECT 17.090 111.920 17.260 113.330 ;
        RECT 14.310 111.800 17.260 111.920 ;
        RECT 14.430 111.750 17.260 111.800 ;
        RECT 17.820 113.420 20.560 113.490 ;
        RECT 21.140 113.420 23.880 113.490 ;
        RECT 17.820 113.320 20.690 113.420 ;
        RECT 17.820 111.910 17.990 113.320 ;
        RECT 18.330 112.450 18.500 112.780 ;
        RECT 18.670 112.750 19.710 112.920 ;
        RECT 18.670 112.310 19.710 112.480 ;
        RECT 19.880 112.450 20.050 112.780 ;
        RECT 20.390 111.910 20.690 113.320 ;
        RECT 17.820 111.770 20.690 111.910 ;
        RECT 21.010 113.320 23.880 113.420 ;
        RECT 21.010 111.910 21.310 113.320 ;
        RECT 21.650 112.450 21.820 112.780 ;
        RECT 21.990 112.750 23.030 112.920 ;
        RECT 21.990 112.310 23.030 112.480 ;
        RECT 23.200 112.450 23.370 112.780 ;
        RECT 23.710 111.910 23.880 113.320 ;
        RECT 21.010 111.770 23.880 111.910 ;
        RECT 17.820 111.740 20.560 111.770 ;
        RECT 21.140 111.740 23.880 111.770 ;
        RECT 24.440 113.450 27.270 113.500 ;
        RECT 24.440 113.330 27.390 113.450 ;
        RECT 24.440 111.920 24.610 113.330 ;
        RECT 24.950 112.460 25.120 112.790 ;
        RECT 25.335 112.760 26.375 112.930 ;
        RECT 25.335 112.320 26.375 112.490 ;
        RECT 26.590 112.460 26.760 112.790 ;
        RECT 27.100 111.920 27.390 113.330 ;
        RECT 24.440 111.800 27.390 111.920 ;
        RECT 24.440 111.750 27.270 111.800 ;
        RECT 14.430 111.350 17.260 111.400 ;
        RECT 14.310 111.230 17.260 111.350 ;
        RECT 14.310 109.820 14.600 111.230 ;
        RECT 14.940 110.360 15.110 110.690 ;
        RECT 15.325 110.660 16.365 110.830 ;
        RECT 15.325 110.220 16.365 110.390 ;
        RECT 16.580 110.360 16.750 110.690 ;
        RECT 17.090 109.820 17.260 111.230 ;
        RECT 14.310 109.700 17.260 109.820 ;
        RECT 14.430 109.650 17.260 109.700 ;
        RECT 17.820 111.320 20.560 111.390 ;
        RECT 21.140 111.320 23.880 111.390 ;
        RECT 17.820 111.220 20.690 111.320 ;
        RECT 17.820 109.810 17.990 111.220 ;
        RECT 18.330 110.350 18.500 110.680 ;
        RECT 18.670 110.650 19.710 110.820 ;
        RECT 18.670 110.210 19.710 110.380 ;
        RECT 19.880 110.350 20.050 110.680 ;
        RECT 20.390 109.810 20.690 111.220 ;
        RECT 17.820 109.670 20.690 109.810 ;
        RECT 21.010 111.220 23.880 111.320 ;
        RECT 21.010 109.810 21.310 111.220 ;
        RECT 21.650 110.350 21.820 110.680 ;
        RECT 21.990 110.650 23.030 110.820 ;
        RECT 21.990 110.210 23.030 110.380 ;
        RECT 23.200 110.350 23.370 110.680 ;
        RECT 23.710 109.810 23.880 111.220 ;
        RECT 21.010 109.670 23.880 109.810 ;
        RECT 17.820 109.640 20.560 109.670 ;
        RECT 21.140 109.640 23.880 109.670 ;
        RECT 24.440 111.350 27.270 111.400 ;
        RECT 24.440 111.230 27.390 111.350 ;
        RECT 24.440 109.820 24.610 111.230 ;
        RECT 24.950 110.360 25.120 110.690 ;
        RECT 25.335 110.660 26.375 110.830 ;
        RECT 25.335 110.220 26.375 110.390 ;
        RECT 26.590 110.360 26.760 110.690 ;
        RECT 27.100 109.820 27.390 111.230 ;
        RECT 24.440 109.700 27.390 109.820 ;
        RECT 24.440 109.650 27.270 109.700 ;
        RECT 14.430 109.250 17.260 109.300 ;
        RECT 14.310 109.130 17.260 109.250 ;
        RECT 14.310 107.720 14.600 109.130 ;
        RECT 14.940 108.260 15.110 108.590 ;
        RECT 15.325 108.560 16.365 108.730 ;
        RECT 15.325 108.120 16.365 108.290 ;
        RECT 16.580 108.260 16.750 108.590 ;
        RECT 17.090 107.720 17.260 109.130 ;
        RECT 14.310 107.600 17.260 107.720 ;
        RECT 14.430 107.550 17.260 107.600 ;
        RECT 17.820 109.220 20.560 109.290 ;
        RECT 21.140 109.220 23.880 109.290 ;
        RECT 17.820 109.120 20.690 109.220 ;
        RECT 17.820 107.710 17.990 109.120 ;
        RECT 18.330 108.250 18.500 108.580 ;
        RECT 18.670 108.550 19.710 108.720 ;
        RECT 18.670 108.110 19.710 108.280 ;
        RECT 19.880 108.250 20.050 108.580 ;
        RECT 20.390 107.710 20.690 109.120 ;
        RECT 17.820 107.570 20.690 107.710 ;
        RECT 21.010 109.120 23.880 109.220 ;
        RECT 21.010 107.710 21.310 109.120 ;
        RECT 21.650 108.250 21.820 108.580 ;
        RECT 21.990 108.550 23.030 108.720 ;
        RECT 21.990 108.110 23.030 108.280 ;
        RECT 23.200 108.250 23.370 108.580 ;
        RECT 23.710 107.710 23.880 109.120 ;
        RECT 21.010 107.570 23.880 107.710 ;
        RECT 17.820 107.540 20.560 107.570 ;
        RECT 21.140 107.540 23.880 107.570 ;
        RECT 24.440 109.250 27.270 109.300 ;
        RECT 24.440 109.130 27.390 109.250 ;
        RECT 24.440 107.720 24.610 109.130 ;
        RECT 24.950 108.260 25.120 108.590 ;
        RECT 25.335 108.560 26.375 108.730 ;
        RECT 25.335 108.120 26.375 108.290 ;
        RECT 26.590 108.260 26.760 108.590 ;
        RECT 27.100 107.720 27.390 109.130 ;
        RECT 24.440 107.600 27.390 107.720 ;
        RECT 24.440 107.550 27.270 107.600 ;
        RECT 14.430 107.150 17.260 107.200 ;
        RECT 14.310 107.030 17.260 107.150 ;
        RECT 14.310 105.620 14.600 107.030 ;
        RECT 14.940 106.160 15.110 106.490 ;
        RECT 15.325 106.460 16.365 106.630 ;
        RECT 15.325 106.020 16.365 106.190 ;
        RECT 16.580 106.160 16.750 106.490 ;
        RECT 17.090 105.620 17.260 107.030 ;
        RECT 14.310 105.500 17.260 105.620 ;
        RECT 14.430 105.450 17.260 105.500 ;
        RECT 17.820 107.120 20.560 107.190 ;
        RECT 21.140 107.120 23.880 107.190 ;
        RECT 17.820 107.020 20.690 107.120 ;
        RECT 17.820 105.610 17.990 107.020 ;
        RECT 18.330 106.150 18.500 106.480 ;
        RECT 18.670 106.450 19.710 106.620 ;
        RECT 18.670 106.010 19.710 106.180 ;
        RECT 19.880 106.150 20.050 106.480 ;
        RECT 20.390 105.610 20.690 107.020 ;
        RECT 17.820 105.470 20.690 105.610 ;
        RECT 21.010 107.020 23.880 107.120 ;
        RECT 21.010 105.610 21.310 107.020 ;
        RECT 21.650 106.150 21.820 106.480 ;
        RECT 21.990 106.450 23.030 106.620 ;
        RECT 21.990 106.010 23.030 106.180 ;
        RECT 23.200 106.150 23.370 106.480 ;
        RECT 23.710 105.610 23.880 107.020 ;
        RECT 21.010 105.470 23.880 105.610 ;
        RECT 17.820 105.440 20.560 105.470 ;
        RECT 21.140 105.440 23.880 105.470 ;
        RECT 24.440 107.150 27.270 107.200 ;
        RECT 24.440 107.030 27.390 107.150 ;
        RECT 24.440 105.620 24.610 107.030 ;
        RECT 24.950 106.160 25.120 106.490 ;
        RECT 25.335 106.460 26.375 106.630 ;
        RECT 25.335 106.020 26.375 106.190 ;
        RECT 26.590 106.160 26.760 106.490 ;
        RECT 27.100 105.620 27.390 107.030 ;
        RECT 24.440 105.500 27.390 105.620 ;
        RECT 24.440 105.450 27.270 105.500 ;
        RECT 14.430 105.050 17.260 105.100 ;
        RECT 14.310 104.930 17.260 105.050 ;
        RECT 14.310 103.520 14.600 104.930 ;
        RECT 14.940 104.060 15.110 104.390 ;
        RECT 15.325 104.360 16.365 104.530 ;
        RECT 15.325 103.920 16.365 104.090 ;
        RECT 16.580 104.060 16.750 104.390 ;
        RECT 17.090 103.520 17.260 104.930 ;
        RECT 14.310 103.400 17.260 103.520 ;
        RECT 14.430 103.350 17.260 103.400 ;
        RECT 17.820 105.020 20.560 105.090 ;
        RECT 21.140 105.020 23.880 105.090 ;
        RECT 17.820 104.920 20.690 105.020 ;
        RECT 17.820 103.510 17.990 104.920 ;
        RECT 18.330 104.050 18.500 104.380 ;
        RECT 18.670 104.350 19.710 104.520 ;
        RECT 18.670 103.910 19.710 104.080 ;
        RECT 19.880 104.050 20.050 104.380 ;
        RECT 20.390 103.510 20.690 104.920 ;
        RECT 17.820 103.370 20.690 103.510 ;
        RECT 21.010 104.920 23.880 105.020 ;
        RECT 21.010 103.510 21.310 104.920 ;
        RECT 21.650 104.050 21.820 104.380 ;
        RECT 21.990 104.350 23.030 104.520 ;
        RECT 21.990 103.910 23.030 104.080 ;
        RECT 23.200 104.050 23.370 104.380 ;
        RECT 23.710 103.510 23.880 104.920 ;
        RECT 21.010 103.370 23.880 103.510 ;
        RECT 17.820 103.340 20.560 103.370 ;
        RECT 21.140 103.340 23.880 103.370 ;
        RECT 24.440 105.050 27.270 105.100 ;
        RECT 24.440 104.930 27.390 105.050 ;
        RECT 24.440 103.520 24.610 104.930 ;
        RECT 24.950 104.060 25.120 104.390 ;
        RECT 25.335 104.360 26.375 104.530 ;
        RECT 25.335 103.920 26.375 104.090 ;
        RECT 26.590 104.060 26.760 104.390 ;
        RECT 27.100 103.520 27.390 104.930 ;
        RECT 24.440 103.400 27.390 103.520 ;
        RECT 24.440 103.350 27.270 103.400 ;
        RECT 14.430 102.950 17.260 103.000 ;
        RECT 14.310 102.830 17.260 102.950 ;
        RECT 14.310 101.420 14.600 102.830 ;
        RECT 14.940 101.960 15.110 102.290 ;
        RECT 15.325 102.260 16.365 102.430 ;
        RECT 15.325 101.820 16.365 101.990 ;
        RECT 16.580 101.960 16.750 102.290 ;
        RECT 17.090 101.420 17.260 102.830 ;
        RECT 14.310 101.300 17.260 101.420 ;
        RECT 14.430 101.250 17.260 101.300 ;
        RECT 17.820 102.920 20.560 102.990 ;
        RECT 21.140 102.920 23.880 102.990 ;
        RECT 17.820 102.820 20.690 102.920 ;
        RECT 17.820 101.410 17.990 102.820 ;
        RECT 18.330 101.950 18.500 102.280 ;
        RECT 18.670 102.250 19.710 102.420 ;
        RECT 18.670 101.810 19.710 101.980 ;
        RECT 19.880 101.950 20.050 102.280 ;
        RECT 20.390 101.410 20.690 102.820 ;
        RECT 17.820 101.270 20.690 101.410 ;
        RECT 21.010 102.820 23.880 102.920 ;
        RECT 21.010 101.410 21.310 102.820 ;
        RECT 21.650 101.950 21.820 102.280 ;
        RECT 21.990 102.250 23.030 102.420 ;
        RECT 21.990 101.810 23.030 101.980 ;
        RECT 23.200 101.950 23.370 102.280 ;
        RECT 23.710 101.410 23.880 102.820 ;
        RECT 21.010 101.270 23.880 101.410 ;
        RECT 17.820 101.240 20.560 101.270 ;
        RECT 21.140 101.240 23.880 101.270 ;
        RECT 24.440 102.950 27.270 103.000 ;
        RECT 24.440 102.830 27.390 102.950 ;
        RECT 24.440 101.420 24.610 102.830 ;
        RECT 24.950 101.960 25.120 102.290 ;
        RECT 25.335 102.260 26.375 102.430 ;
        RECT 25.335 101.820 26.375 101.990 ;
        RECT 26.590 101.960 26.760 102.290 ;
        RECT 27.100 101.420 27.390 102.830 ;
        RECT 24.440 101.300 27.390 101.420 ;
        RECT 24.440 101.250 27.270 101.300 ;
        RECT 14.430 100.850 17.260 100.900 ;
        RECT 14.310 100.730 17.260 100.850 ;
        RECT 14.310 99.320 14.600 100.730 ;
        RECT 14.940 99.860 15.110 100.190 ;
        RECT 15.325 100.160 16.365 100.330 ;
        RECT 15.325 99.720 16.365 99.890 ;
        RECT 16.580 99.860 16.750 100.190 ;
        RECT 17.090 99.320 17.260 100.730 ;
        RECT 14.310 99.200 17.260 99.320 ;
        RECT 14.430 99.150 17.260 99.200 ;
        RECT 17.820 100.820 20.560 100.890 ;
        RECT 21.140 100.820 23.880 100.890 ;
        RECT 17.820 100.720 20.690 100.820 ;
        RECT 17.820 99.310 17.990 100.720 ;
        RECT 18.330 99.850 18.500 100.180 ;
        RECT 18.670 100.150 19.710 100.320 ;
        RECT 18.670 99.710 19.710 99.880 ;
        RECT 19.880 99.850 20.050 100.180 ;
        RECT 20.390 99.310 20.690 100.720 ;
        RECT 17.820 99.170 20.690 99.310 ;
        RECT 21.010 100.720 23.880 100.820 ;
        RECT 21.010 99.310 21.310 100.720 ;
        RECT 21.650 99.850 21.820 100.180 ;
        RECT 21.990 100.150 23.030 100.320 ;
        RECT 21.990 99.710 23.030 99.880 ;
        RECT 23.200 99.850 23.370 100.180 ;
        RECT 23.710 99.310 23.880 100.720 ;
        RECT 21.010 99.170 23.880 99.310 ;
        RECT 17.820 99.140 20.560 99.170 ;
        RECT 21.140 99.140 23.880 99.170 ;
        RECT 24.440 100.850 27.270 100.900 ;
        RECT 24.440 100.730 27.390 100.850 ;
        RECT 24.440 99.320 24.610 100.730 ;
        RECT 24.950 99.860 25.120 100.190 ;
        RECT 25.335 100.160 26.375 100.330 ;
        RECT 25.335 99.720 26.375 99.890 ;
        RECT 26.590 99.860 26.760 100.190 ;
        RECT 27.100 99.320 27.390 100.730 ;
        RECT 24.440 99.200 27.390 99.320 ;
        RECT 24.440 99.150 27.270 99.200 ;
        RECT 14.430 98.750 17.260 98.800 ;
        RECT 14.310 98.630 17.260 98.750 ;
        RECT 14.310 97.220 14.600 98.630 ;
        RECT 14.940 97.760 15.110 98.090 ;
        RECT 15.325 98.060 16.365 98.230 ;
        RECT 15.325 97.620 16.365 97.790 ;
        RECT 16.580 97.760 16.750 98.090 ;
        RECT 17.090 97.220 17.260 98.630 ;
        RECT 14.310 97.100 17.260 97.220 ;
        RECT 14.430 97.050 17.260 97.100 ;
        RECT 17.820 98.720 20.560 98.790 ;
        RECT 21.140 98.720 23.880 98.790 ;
        RECT 17.820 98.620 20.690 98.720 ;
        RECT 17.820 97.210 17.990 98.620 ;
        RECT 18.330 97.750 18.500 98.080 ;
        RECT 18.670 98.050 19.710 98.220 ;
        RECT 18.670 97.610 19.710 97.780 ;
        RECT 19.880 97.750 20.050 98.080 ;
        RECT 20.390 97.210 20.690 98.620 ;
        RECT 17.820 97.070 20.690 97.210 ;
        RECT 21.010 98.620 23.880 98.720 ;
        RECT 21.010 97.210 21.310 98.620 ;
        RECT 21.650 97.750 21.820 98.080 ;
        RECT 21.990 98.050 23.030 98.220 ;
        RECT 21.990 97.610 23.030 97.780 ;
        RECT 23.200 97.750 23.370 98.080 ;
        RECT 23.710 97.210 23.880 98.620 ;
        RECT 21.010 97.070 23.880 97.210 ;
        RECT 17.820 97.040 20.560 97.070 ;
        RECT 21.140 97.040 23.880 97.070 ;
        RECT 24.440 98.750 27.270 98.800 ;
        RECT 24.440 98.630 27.390 98.750 ;
        RECT 24.440 97.220 24.610 98.630 ;
        RECT 24.950 97.760 25.120 98.090 ;
        RECT 25.335 98.060 26.375 98.230 ;
        RECT 25.335 97.620 26.375 97.790 ;
        RECT 26.590 97.760 26.760 98.090 ;
        RECT 27.100 97.220 27.390 98.630 ;
        RECT 24.440 97.100 27.390 97.220 ;
        RECT 24.440 97.050 27.270 97.100 ;
        RECT 14.430 96.650 17.260 96.700 ;
        RECT 14.310 96.530 17.260 96.650 ;
        RECT 14.310 95.120 14.600 96.530 ;
        RECT 14.940 95.660 15.110 95.990 ;
        RECT 15.325 95.960 16.365 96.130 ;
        RECT 15.325 95.520 16.365 95.690 ;
        RECT 16.580 95.660 16.750 95.990 ;
        RECT 17.090 95.120 17.260 96.530 ;
        RECT 14.310 95.000 17.260 95.120 ;
        RECT 14.430 94.950 17.260 95.000 ;
        RECT 17.820 96.620 20.560 96.690 ;
        RECT 21.140 96.620 23.880 96.690 ;
        RECT 17.820 96.520 20.690 96.620 ;
        RECT 17.820 95.110 17.990 96.520 ;
        RECT 18.330 95.650 18.500 95.980 ;
        RECT 18.670 95.950 19.710 96.120 ;
        RECT 18.670 95.510 19.710 95.680 ;
        RECT 19.880 95.650 20.050 95.980 ;
        RECT 20.390 95.110 20.690 96.520 ;
        RECT 17.820 94.970 20.690 95.110 ;
        RECT 21.010 96.520 23.880 96.620 ;
        RECT 21.010 95.110 21.310 96.520 ;
        RECT 21.650 95.650 21.820 95.980 ;
        RECT 21.990 95.950 23.030 96.120 ;
        RECT 21.990 95.510 23.030 95.680 ;
        RECT 23.200 95.650 23.370 95.980 ;
        RECT 23.710 95.110 23.880 96.520 ;
        RECT 21.010 94.970 23.880 95.110 ;
        RECT 17.820 94.940 20.560 94.970 ;
        RECT 21.140 94.940 23.880 94.970 ;
        RECT 24.440 96.650 27.270 96.700 ;
        RECT 24.440 96.530 27.390 96.650 ;
        RECT 24.440 95.120 24.610 96.530 ;
        RECT 24.950 95.660 25.120 95.990 ;
        RECT 25.335 95.960 26.375 96.130 ;
        RECT 25.335 95.520 26.375 95.690 ;
        RECT 26.590 95.660 26.760 95.990 ;
        RECT 27.100 95.120 27.390 96.530 ;
        RECT 24.440 95.000 27.390 95.120 ;
        RECT 24.440 94.950 27.270 95.000 ;
        RECT 14.430 94.550 17.260 94.600 ;
        RECT 14.310 94.430 17.260 94.550 ;
        RECT 14.310 93.020 14.600 94.430 ;
        RECT 14.940 93.560 15.110 93.890 ;
        RECT 15.325 93.860 16.365 94.030 ;
        RECT 15.325 93.420 16.365 93.590 ;
        RECT 16.580 93.560 16.750 93.890 ;
        RECT 17.090 93.020 17.260 94.430 ;
        RECT 14.310 92.900 17.260 93.020 ;
        RECT 14.430 92.850 17.260 92.900 ;
        RECT 17.820 94.520 20.560 94.590 ;
        RECT 21.140 94.520 23.880 94.590 ;
        RECT 17.820 94.420 20.690 94.520 ;
        RECT 17.820 93.010 17.990 94.420 ;
        RECT 18.330 93.550 18.500 93.880 ;
        RECT 18.670 93.850 19.710 94.020 ;
        RECT 18.670 93.410 19.710 93.580 ;
        RECT 19.880 93.550 20.050 93.880 ;
        RECT 20.390 93.010 20.690 94.420 ;
        RECT 17.820 92.870 20.690 93.010 ;
        RECT 21.010 94.420 23.880 94.520 ;
        RECT 21.010 93.010 21.310 94.420 ;
        RECT 21.650 93.550 21.820 93.880 ;
        RECT 21.990 93.850 23.030 94.020 ;
        RECT 21.990 93.410 23.030 93.580 ;
        RECT 23.200 93.550 23.370 93.880 ;
        RECT 23.710 93.010 23.880 94.420 ;
        RECT 21.010 92.870 23.880 93.010 ;
        RECT 17.820 92.840 20.560 92.870 ;
        RECT 21.140 92.840 23.880 92.870 ;
        RECT 24.440 94.550 27.270 94.600 ;
        RECT 24.440 94.430 27.390 94.550 ;
        RECT 24.440 93.020 24.610 94.430 ;
        RECT 24.950 93.560 25.120 93.890 ;
        RECT 25.335 93.860 26.375 94.030 ;
        RECT 25.335 93.420 26.375 93.590 ;
        RECT 26.590 93.560 26.760 93.890 ;
        RECT 27.100 93.020 27.390 94.430 ;
        RECT 24.440 92.900 27.390 93.020 ;
        RECT 24.440 92.850 27.270 92.900 ;
        RECT 14.430 92.450 17.260 92.500 ;
        RECT 14.310 92.330 17.260 92.450 ;
        RECT 14.310 90.920 14.600 92.330 ;
        RECT 14.940 91.460 15.110 91.790 ;
        RECT 15.325 91.760 16.365 91.930 ;
        RECT 15.325 91.320 16.365 91.490 ;
        RECT 16.580 91.460 16.750 91.790 ;
        RECT 17.090 90.920 17.260 92.330 ;
        RECT 14.310 90.800 17.260 90.920 ;
        RECT 14.430 90.750 17.260 90.800 ;
        RECT 17.820 92.420 20.560 92.490 ;
        RECT 21.140 92.420 23.880 92.490 ;
        RECT 17.820 92.320 20.690 92.420 ;
        RECT 17.820 90.910 17.990 92.320 ;
        RECT 18.330 91.450 18.500 91.780 ;
        RECT 18.670 91.750 19.710 91.920 ;
        RECT 18.670 91.310 19.710 91.480 ;
        RECT 19.880 91.450 20.050 91.780 ;
        RECT 20.390 90.910 20.690 92.320 ;
        RECT 17.820 90.770 20.690 90.910 ;
        RECT 21.010 92.320 23.880 92.420 ;
        RECT 21.010 90.910 21.310 92.320 ;
        RECT 21.650 91.450 21.820 91.780 ;
        RECT 21.990 91.750 23.030 91.920 ;
        RECT 21.990 91.310 23.030 91.480 ;
        RECT 23.200 91.450 23.370 91.780 ;
        RECT 23.710 90.910 23.880 92.320 ;
        RECT 21.010 90.770 23.880 90.910 ;
        RECT 17.820 90.740 20.560 90.770 ;
        RECT 21.140 90.740 23.880 90.770 ;
        RECT 24.440 92.450 27.270 92.500 ;
        RECT 24.440 92.330 27.390 92.450 ;
        RECT 24.440 90.920 24.610 92.330 ;
        RECT 24.950 91.460 25.120 91.790 ;
        RECT 25.335 91.760 26.375 91.930 ;
        RECT 25.335 91.320 26.375 91.490 ;
        RECT 26.590 91.460 26.760 91.790 ;
        RECT 27.100 90.920 27.390 92.330 ;
        RECT 24.440 90.800 27.390 90.920 ;
        RECT 24.440 90.750 27.270 90.800 ;
        RECT 14.430 90.350 17.260 90.400 ;
        RECT 14.310 90.230 17.260 90.350 ;
        RECT 14.310 88.820 14.600 90.230 ;
        RECT 14.940 89.360 15.110 89.690 ;
        RECT 15.325 89.660 16.365 89.830 ;
        RECT 15.325 89.220 16.365 89.390 ;
        RECT 16.580 89.360 16.750 89.690 ;
        RECT 17.090 88.820 17.260 90.230 ;
        RECT 14.310 88.700 17.260 88.820 ;
        RECT 14.430 88.650 17.260 88.700 ;
        RECT 17.820 90.320 20.560 90.390 ;
        RECT 21.140 90.320 23.880 90.390 ;
        RECT 17.820 90.220 20.690 90.320 ;
        RECT 17.820 88.810 17.990 90.220 ;
        RECT 18.330 89.350 18.500 89.680 ;
        RECT 18.670 89.650 19.710 89.820 ;
        RECT 18.670 89.210 19.710 89.380 ;
        RECT 19.880 89.350 20.050 89.680 ;
        RECT 20.390 88.810 20.690 90.220 ;
        RECT 17.820 88.670 20.690 88.810 ;
        RECT 21.010 90.220 23.880 90.320 ;
        RECT 21.010 88.810 21.310 90.220 ;
        RECT 21.650 89.350 21.820 89.680 ;
        RECT 21.990 89.650 23.030 89.820 ;
        RECT 21.990 89.210 23.030 89.380 ;
        RECT 23.200 89.350 23.370 89.680 ;
        RECT 23.710 88.810 23.880 90.220 ;
        RECT 21.010 88.670 23.880 88.810 ;
        RECT 17.820 88.640 20.560 88.670 ;
        RECT 21.140 88.640 23.880 88.670 ;
        RECT 24.440 90.350 27.270 90.400 ;
        RECT 24.440 90.230 27.390 90.350 ;
        RECT 24.440 88.820 24.610 90.230 ;
        RECT 24.950 89.360 25.120 89.690 ;
        RECT 25.335 89.660 26.375 89.830 ;
        RECT 25.335 89.220 26.375 89.390 ;
        RECT 26.590 89.360 26.760 89.690 ;
        RECT 27.100 88.820 27.390 90.230 ;
        RECT 24.440 88.700 27.390 88.820 ;
        RECT 24.440 88.650 27.270 88.700 ;
        RECT 14.430 88.250 17.260 88.300 ;
        RECT 14.310 88.130 17.260 88.250 ;
        RECT 14.310 86.720 14.600 88.130 ;
        RECT 14.940 87.260 15.110 87.590 ;
        RECT 15.325 87.560 16.365 87.730 ;
        RECT 15.325 87.120 16.365 87.290 ;
        RECT 16.580 87.260 16.750 87.590 ;
        RECT 17.090 86.720 17.260 88.130 ;
        RECT 14.310 86.600 17.260 86.720 ;
        RECT 14.430 86.550 17.260 86.600 ;
        RECT 17.820 88.220 20.560 88.290 ;
        RECT 21.140 88.220 23.880 88.290 ;
        RECT 17.820 88.120 20.690 88.220 ;
        RECT 17.820 86.710 17.990 88.120 ;
        RECT 18.330 87.250 18.500 87.580 ;
        RECT 18.670 87.550 19.710 87.720 ;
        RECT 18.670 87.110 19.710 87.280 ;
        RECT 19.880 87.250 20.050 87.580 ;
        RECT 20.390 86.710 20.690 88.120 ;
        RECT 17.820 86.570 20.690 86.710 ;
        RECT 21.010 88.120 23.880 88.220 ;
        RECT 21.010 86.710 21.310 88.120 ;
        RECT 21.650 87.250 21.820 87.580 ;
        RECT 21.990 87.550 23.030 87.720 ;
        RECT 21.990 87.110 23.030 87.280 ;
        RECT 23.200 87.250 23.370 87.580 ;
        RECT 23.710 86.710 23.880 88.120 ;
        RECT 21.010 86.570 23.880 86.710 ;
        RECT 17.820 86.540 20.560 86.570 ;
        RECT 21.140 86.540 23.880 86.570 ;
        RECT 24.440 88.250 27.270 88.300 ;
        RECT 24.440 88.130 27.390 88.250 ;
        RECT 24.440 86.720 24.610 88.130 ;
        RECT 24.950 87.260 25.120 87.590 ;
        RECT 25.335 87.560 26.375 87.730 ;
        RECT 25.335 87.120 26.375 87.290 ;
        RECT 26.590 87.260 26.760 87.590 ;
        RECT 27.100 86.720 27.390 88.130 ;
        RECT 24.440 86.600 27.390 86.720 ;
        RECT 24.440 86.550 27.270 86.600 ;
        RECT 14.430 86.150 17.260 86.200 ;
        RECT 14.310 86.030 17.260 86.150 ;
        RECT 14.310 84.620 14.600 86.030 ;
        RECT 14.940 85.160 15.110 85.490 ;
        RECT 15.325 85.460 16.365 85.630 ;
        RECT 15.325 85.020 16.365 85.190 ;
        RECT 16.580 85.160 16.750 85.490 ;
        RECT 17.090 84.620 17.260 86.030 ;
        RECT 14.310 84.500 17.260 84.620 ;
        RECT 14.430 84.450 17.260 84.500 ;
        RECT 17.820 86.120 20.560 86.190 ;
        RECT 21.140 86.120 23.880 86.190 ;
        RECT 17.820 86.020 20.690 86.120 ;
        RECT 17.820 84.610 17.990 86.020 ;
        RECT 18.330 85.150 18.500 85.480 ;
        RECT 18.670 85.450 19.710 85.620 ;
        RECT 18.670 85.010 19.710 85.180 ;
        RECT 19.880 85.150 20.050 85.480 ;
        RECT 20.390 84.610 20.690 86.020 ;
        RECT 17.820 84.470 20.690 84.610 ;
        RECT 21.010 86.020 23.880 86.120 ;
        RECT 21.010 84.610 21.310 86.020 ;
        RECT 21.650 85.150 21.820 85.480 ;
        RECT 21.990 85.450 23.030 85.620 ;
        RECT 21.990 85.010 23.030 85.180 ;
        RECT 23.200 85.150 23.370 85.480 ;
        RECT 23.710 84.610 23.880 86.020 ;
        RECT 21.010 84.470 23.880 84.610 ;
        RECT 17.820 84.440 20.560 84.470 ;
        RECT 21.140 84.440 23.880 84.470 ;
        RECT 24.440 86.150 27.270 86.200 ;
        RECT 24.440 86.030 27.390 86.150 ;
        RECT 24.440 84.620 24.610 86.030 ;
        RECT 24.950 85.160 25.120 85.490 ;
        RECT 25.335 85.460 26.375 85.630 ;
        RECT 25.335 85.020 26.375 85.190 ;
        RECT 26.590 85.160 26.760 85.490 ;
        RECT 27.100 84.620 27.390 86.030 ;
        RECT 24.440 84.500 27.390 84.620 ;
        RECT 24.440 84.450 27.270 84.500 ;
        RECT 14.430 84.050 17.260 84.100 ;
        RECT 14.310 83.930 17.260 84.050 ;
        RECT 14.310 82.520 14.600 83.930 ;
        RECT 14.940 83.060 15.110 83.390 ;
        RECT 15.325 83.360 16.365 83.530 ;
        RECT 15.325 82.920 16.365 83.090 ;
        RECT 16.580 83.060 16.750 83.390 ;
        RECT 17.090 82.520 17.260 83.930 ;
        RECT 14.310 82.400 17.260 82.520 ;
        RECT 14.430 82.350 17.260 82.400 ;
        RECT 17.820 84.020 20.560 84.090 ;
        RECT 21.140 84.020 23.880 84.090 ;
        RECT 17.820 83.920 20.690 84.020 ;
        RECT 17.820 82.510 17.990 83.920 ;
        RECT 18.330 83.050 18.500 83.380 ;
        RECT 18.670 83.350 19.710 83.520 ;
        RECT 18.670 82.910 19.710 83.080 ;
        RECT 19.880 83.050 20.050 83.380 ;
        RECT 20.390 82.510 20.690 83.920 ;
        RECT 17.820 82.370 20.690 82.510 ;
        RECT 21.010 83.920 23.880 84.020 ;
        RECT 21.010 82.510 21.310 83.920 ;
        RECT 21.650 83.050 21.820 83.380 ;
        RECT 21.990 83.350 23.030 83.520 ;
        RECT 21.990 82.910 23.030 83.080 ;
        RECT 23.200 83.050 23.370 83.380 ;
        RECT 23.710 82.510 23.880 83.920 ;
        RECT 21.010 82.370 23.880 82.510 ;
        RECT 17.820 82.340 20.560 82.370 ;
        RECT 21.140 82.340 23.880 82.370 ;
        RECT 24.440 84.050 27.270 84.100 ;
        RECT 24.440 83.930 27.390 84.050 ;
        RECT 24.440 82.520 24.610 83.930 ;
        RECT 24.950 83.060 25.120 83.390 ;
        RECT 25.335 83.360 26.375 83.530 ;
        RECT 25.335 82.920 26.375 83.090 ;
        RECT 26.590 83.060 26.760 83.390 ;
        RECT 27.100 82.520 27.390 83.930 ;
        RECT 24.440 82.400 27.390 82.520 ;
        RECT 24.440 82.350 27.270 82.400 ;
        RECT 14.430 81.950 17.260 82.000 ;
        RECT 14.310 81.830 17.260 81.950 ;
        RECT 14.310 80.420 14.600 81.830 ;
        RECT 14.940 80.960 15.110 81.290 ;
        RECT 15.325 81.260 16.365 81.430 ;
        RECT 15.325 80.820 16.365 80.990 ;
        RECT 16.580 80.960 16.750 81.290 ;
        RECT 17.090 80.420 17.260 81.830 ;
        RECT 14.310 80.300 17.260 80.420 ;
        RECT 14.430 80.250 17.260 80.300 ;
        RECT 17.820 81.920 20.560 81.990 ;
        RECT 21.140 81.920 23.880 81.990 ;
        RECT 17.820 81.820 20.690 81.920 ;
        RECT 17.820 80.410 17.990 81.820 ;
        RECT 18.330 80.950 18.500 81.280 ;
        RECT 18.670 81.250 19.710 81.420 ;
        RECT 18.670 80.810 19.710 80.980 ;
        RECT 19.880 80.950 20.050 81.280 ;
        RECT 20.390 80.410 20.690 81.820 ;
        RECT 17.820 80.270 20.690 80.410 ;
        RECT 21.010 81.820 23.880 81.920 ;
        RECT 21.010 80.410 21.310 81.820 ;
        RECT 21.650 80.950 21.820 81.280 ;
        RECT 21.990 81.250 23.030 81.420 ;
        RECT 21.990 80.810 23.030 80.980 ;
        RECT 23.200 80.950 23.370 81.280 ;
        RECT 23.710 80.410 23.880 81.820 ;
        RECT 21.010 80.270 23.880 80.410 ;
        RECT 17.820 80.240 20.560 80.270 ;
        RECT 21.140 80.240 23.880 80.270 ;
        RECT 24.440 81.950 27.270 82.000 ;
        RECT 24.440 81.830 27.390 81.950 ;
        RECT 24.440 80.420 24.610 81.830 ;
        RECT 24.950 80.960 25.120 81.290 ;
        RECT 25.335 81.260 26.375 81.430 ;
        RECT 25.335 80.820 26.375 80.990 ;
        RECT 26.590 80.960 26.760 81.290 ;
        RECT 27.100 80.420 27.390 81.830 ;
        RECT 24.440 80.300 27.390 80.420 ;
        RECT 24.440 80.250 27.270 80.300 ;
        RECT 14.430 79.850 17.260 79.900 ;
        RECT 14.310 79.730 17.260 79.850 ;
        RECT 14.310 78.320 14.600 79.730 ;
        RECT 14.940 78.860 15.110 79.190 ;
        RECT 15.325 79.160 16.365 79.330 ;
        RECT 15.325 78.720 16.365 78.890 ;
        RECT 16.580 78.860 16.750 79.190 ;
        RECT 17.090 78.320 17.260 79.730 ;
        RECT 14.310 78.200 17.260 78.320 ;
        RECT 14.430 78.150 17.260 78.200 ;
        RECT 17.820 79.820 20.560 79.890 ;
        RECT 21.140 79.820 23.880 79.890 ;
        RECT 17.820 79.720 20.690 79.820 ;
        RECT 17.820 78.310 17.990 79.720 ;
        RECT 18.330 78.850 18.500 79.180 ;
        RECT 18.670 79.150 19.710 79.320 ;
        RECT 18.670 78.710 19.710 78.880 ;
        RECT 19.880 78.850 20.050 79.180 ;
        RECT 20.390 78.310 20.690 79.720 ;
        RECT 17.820 78.170 20.690 78.310 ;
        RECT 21.010 79.720 23.880 79.820 ;
        RECT 21.010 78.310 21.310 79.720 ;
        RECT 21.650 78.850 21.820 79.180 ;
        RECT 21.990 79.150 23.030 79.320 ;
        RECT 21.990 78.710 23.030 78.880 ;
        RECT 23.200 78.850 23.370 79.180 ;
        RECT 23.710 78.310 23.880 79.720 ;
        RECT 21.010 78.170 23.880 78.310 ;
        RECT 17.820 78.140 20.560 78.170 ;
        RECT 21.140 78.140 23.880 78.170 ;
        RECT 24.440 79.850 27.270 79.900 ;
        RECT 24.440 79.730 27.390 79.850 ;
        RECT 24.440 78.320 24.610 79.730 ;
        RECT 24.950 78.860 25.120 79.190 ;
        RECT 25.335 79.160 26.375 79.330 ;
        RECT 25.335 78.720 26.375 78.890 ;
        RECT 26.590 78.860 26.760 79.190 ;
        RECT 27.100 78.320 27.390 79.730 ;
        RECT 24.440 78.200 27.390 78.320 ;
        RECT 24.440 78.150 27.270 78.200 ;
        RECT 14.430 77.750 17.260 77.800 ;
        RECT 14.310 77.630 17.260 77.750 ;
        RECT 14.310 76.220 14.600 77.630 ;
        RECT 14.940 76.760 15.110 77.090 ;
        RECT 15.325 77.060 16.365 77.230 ;
        RECT 15.325 76.620 16.365 76.790 ;
        RECT 16.580 76.760 16.750 77.090 ;
        RECT 17.090 76.220 17.260 77.630 ;
        RECT 14.310 76.100 17.260 76.220 ;
        RECT 14.430 76.050 17.260 76.100 ;
        RECT 17.820 77.720 20.560 77.790 ;
        RECT 21.140 77.720 23.880 77.790 ;
        RECT 17.820 77.620 20.690 77.720 ;
        RECT 17.820 76.210 17.990 77.620 ;
        RECT 18.330 76.750 18.500 77.080 ;
        RECT 18.670 77.050 19.710 77.220 ;
        RECT 18.670 76.610 19.710 76.780 ;
        RECT 19.880 76.750 20.050 77.080 ;
        RECT 20.390 76.210 20.690 77.620 ;
        RECT 17.820 76.070 20.690 76.210 ;
        RECT 21.010 77.620 23.880 77.720 ;
        RECT 21.010 76.210 21.310 77.620 ;
        RECT 21.650 76.750 21.820 77.080 ;
        RECT 21.990 77.050 23.030 77.220 ;
        RECT 21.990 76.610 23.030 76.780 ;
        RECT 23.200 76.750 23.370 77.080 ;
        RECT 23.710 76.210 23.880 77.620 ;
        RECT 21.010 76.070 23.880 76.210 ;
        RECT 17.820 76.040 20.560 76.070 ;
        RECT 21.140 76.040 23.880 76.070 ;
        RECT 24.440 77.750 27.270 77.800 ;
        RECT 24.440 77.630 27.390 77.750 ;
        RECT 24.440 76.220 24.610 77.630 ;
        RECT 24.950 76.760 25.120 77.090 ;
        RECT 25.335 77.060 26.375 77.230 ;
        RECT 25.335 76.620 26.375 76.790 ;
        RECT 26.590 76.760 26.760 77.090 ;
        RECT 27.100 76.220 27.390 77.630 ;
        RECT 24.440 76.100 27.390 76.220 ;
        RECT 24.440 76.050 27.270 76.100 ;
        RECT 14.430 75.650 17.260 75.700 ;
        RECT 14.310 75.530 17.260 75.650 ;
        RECT 14.310 74.120 14.600 75.530 ;
        RECT 14.940 74.660 15.110 74.990 ;
        RECT 15.325 74.960 16.365 75.130 ;
        RECT 15.325 74.520 16.365 74.690 ;
        RECT 16.580 74.660 16.750 74.990 ;
        RECT 17.090 74.120 17.260 75.530 ;
        RECT 14.310 74.000 17.260 74.120 ;
        RECT 14.430 73.950 17.260 74.000 ;
        RECT 17.820 75.620 20.560 75.690 ;
        RECT 21.140 75.620 23.880 75.690 ;
        RECT 17.820 75.520 20.690 75.620 ;
        RECT 17.820 74.110 17.990 75.520 ;
        RECT 18.330 74.650 18.500 74.980 ;
        RECT 18.670 74.950 19.710 75.120 ;
        RECT 18.670 74.510 19.710 74.680 ;
        RECT 19.880 74.650 20.050 74.980 ;
        RECT 20.390 74.110 20.690 75.520 ;
        RECT 17.820 73.970 20.690 74.110 ;
        RECT 21.010 75.520 23.880 75.620 ;
        RECT 21.010 74.110 21.310 75.520 ;
        RECT 21.650 74.650 21.820 74.980 ;
        RECT 21.990 74.950 23.030 75.120 ;
        RECT 21.990 74.510 23.030 74.680 ;
        RECT 23.200 74.650 23.370 74.980 ;
        RECT 23.710 74.110 23.880 75.520 ;
        RECT 21.010 73.970 23.880 74.110 ;
        RECT 17.820 73.940 20.560 73.970 ;
        RECT 21.140 73.940 23.880 73.970 ;
        RECT 24.440 75.650 27.270 75.700 ;
        RECT 24.440 75.530 27.390 75.650 ;
        RECT 24.440 74.120 24.610 75.530 ;
        RECT 24.950 74.660 25.120 74.990 ;
        RECT 25.335 74.960 26.375 75.130 ;
        RECT 25.335 74.520 26.375 74.690 ;
        RECT 26.590 74.660 26.760 74.990 ;
        RECT 27.100 74.120 27.390 75.530 ;
        RECT 24.440 74.000 27.390 74.120 ;
        RECT 24.440 73.950 27.270 74.000 ;
        RECT 14.430 73.550 17.260 73.600 ;
        RECT 14.310 73.430 17.260 73.550 ;
        RECT 14.310 72.020 14.600 73.430 ;
        RECT 14.940 72.560 15.110 72.890 ;
        RECT 15.325 72.860 16.365 73.030 ;
        RECT 15.325 72.420 16.365 72.590 ;
        RECT 16.580 72.560 16.750 72.890 ;
        RECT 17.090 72.020 17.260 73.430 ;
        RECT 14.310 71.900 17.260 72.020 ;
        RECT 14.430 71.850 17.260 71.900 ;
        RECT 17.820 73.520 20.560 73.590 ;
        RECT 21.140 73.520 23.880 73.590 ;
        RECT 17.820 73.420 20.690 73.520 ;
        RECT 17.820 72.010 17.990 73.420 ;
        RECT 18.330 72.550 18.500 72.880 ;
        RECT 18.670 72.850 19.710 73.020 ;
        RECT 18.670 72.410 19.710 72.580 ;
        RECT 19.880 72.550 20.050 72.880 ;
        RECT 20.390 72.010 20.690 73.420 ;
        RECT 17.820 71.870 20.690 72.010 ;
        RECT 21.010 73.420 23.880 73.520 ;
        RECT 21.010 72.010 21.310 73.420 ;
        RECT 21.650 72.550 21.820 72.880 ;
        RECT 21.990 72.850 23.030 73.020 ;
        RECT 21.990 72.410 23.030 72.580 ;
        RECT 23.200 72.550 23.370 72.880 ;
        RECT 23.710 72.010 23.880 73.420 ;
        RECT 21.010 71.870 23.880 72.010 ;
        RECT 17.820 71.840 20.560 71.870 ;
        RECT 21.140 71.840 23.880 71.870 ;
        RECT 24.440 73.550 27.270 73.600 ;
        RECT 24.440 73.430 27.390 73.550 ;
        RECT 24.440 72.020 24.610 73.430 ;
        RECT 24.950 72.560 25.120 72.890 ;
        RECT 25.335 72.860 26.375 73.030 ;
        RECT 25.335 72.420 26.375 72.590 ;
        RECT 26.590 72.560 26.760 72.890 ;
        RECT 27.100 72.020 27.390 73.430 ;
        RECT 24.440 71.900 27.390 72.020 ;
        RECT 24.440 71.850 27.270 71.900 ;
        RECT 14.430 71.450 17.260 71.500 ;
        RECT 14.310 71.330 17.260 71.450 ;
        RECT 14.310 69.920 14.600 71.330 ;
        RECT 14.940 70.460 15.110 70.790 ;
        RECT 15.325 70.760 16.365 70.930 ;
        RECT 15.325 70.320 16.365 70.490 ;
        RECT 16.580 70.460 16.750 70.790 ;
        RECT 17.090 69.920 17.260 71.330 ;
        RECT 14.310 69.800 17.260 69.920 ;
        RECT 14.430 69.750 17.260 69.800 ;
        RECT 17.820 71.420 20.560 71.490 ;
        RECT 21.140 71.420 23.880 71.490 ;
        RECT 17.820 71.320 20.690 71.420 ;
        RECT 17.820 69.910 17.990 71.320 ;
        RECT 18.330 70.450 18.500 70.780 ;
        RECT 18.670 70.750 19.710 70.920 ;
        RECT 18.670 70.310 19.710 70.480 ;
        RECT 19.880 70.450 20.050 70.780 ;
        RECT 20.390 69.910 20.690 71.320 ;
        RECT 17.820 69.770 20.690 69.910 ;
        RECT 21.010 71.320 23.880 71.420 ;
        RECT 21.010 69.910 21.310 71.320 ;
        RECT 21.650 70.450 21.820 70.780 ;
        RECT 21.990 70.750 23.030 70.920 ;
        RECT 21.990 70.310 23.030 70.480 ;
        RECT 23.200 70.450 23.370 70.780 ;
        RECT 23.710 69.910 23.880 71.320 ;
        RECT 21.010 69.770 23.880 69.910 ;
        RECT 17.820 69.740 20.560 69.770 ;
        RECT 21.140 69.740 23.880 69.770 ;
        RECT 24.440 71.450 27.270 71.500 ;
        RECT 24.440 71.330 27.390 71.450 ;
        RECT 24.440 69.920 24.610 71.330 ;
        RECT 24.950 70.460 25.120 70.790 ;
        RECT 25.335 70.760 26.375 70.930 ;
        RECT 25.335 70.320 26.375 70.490 ;
        RECT 26.590 70.460 26.760 70.790 ;
        RECT 27.100 69.920 27.390 71.330 ;
        RECT 24.440 69.800 27.390 69.920 ;
        RECT 24.440 69.750 27.270 69.800 ;
        RECT 14.430 69.350 17.260 69.400 ;
        RECT 14.310 69.230 17.260 69.350 ;
        RECT 14.310 67.820 14.600 69.230 ;
        RECT 14.940 68.360 15.110 68.690 ;
        RECT 15.325 68.660 16.365 68.830 ;
        RECT 15.325 68.220 16.365 68.390 ;
        RECT 16.580 68.360 16.750 68.690 ;
        RECT 17.090 67.820 17.260 69.230 ;
        RECT 14.310 67.700 17.260 67.820 ;
        RECT 14.430 67.650 17.260 67.700 ;
        RECT 17.820 69.320 20.560 69.390 ;
        RECT 21.140 69.320 23.880 69.390 ;
        RECT 17.820 69.220 20.690 69.320 ;
        RECT 17.820 67.810 17.990 69.220 ;
        RECT 18.330 68.350 18.500 68.680 ;
        RECT 18.670 68.650 19.710 68.820 ;
        RECT 18.670 68.210 19.710 68.380 ;
        RECT 19.880 68.350 20.050 68.680 ;
        RECT 20.390 67.810 20.690 69.220 ;
        RECT 17.820 67.670 20.690 67.810 ;
        RECT 21.010 69.220 23.880 69.320 ;
        RECT 21.010 67.810 21.310 69.220 ;
        RECT 21.650 68.350 21.820 68.680 ;
        RECT 21.990 68.650 23.030 68.820 ;
        RECT 21.990 68.210 23.030 68.380 ;
        RECT 23.200 68.350 23.370 68.680 ;
        RECT 23.710 67.810 23.880 69.220 ;
        RECT 21.010 67.670 23.880 67.810 ;
        RECT 17.820 67.640 20.560 67.670 ;
        RECT 21.140 67.640 23.880 67.670 ;
        RECT 24.440 69.350 27.270 69.400 ;
        RECT 24.440 69.230 27.390 69.350 ;
        RECT 24.440 67.820 24.610 69.230 ;
        RECT 24.950 68.360 25.120 68.690 ;
        RECT 25.335 68.660 26.375 68.830 ;
        RECT 25.335 68.220 26.375 68.390 ;
        RECT 26.590 68.360 26.760 68.690 ;
        RECT 27.100 67.820 27.390 69.230 ;
        RECT 24.440 67.700 27.390 67.820 ;
        RECT 24.440 67.650 27.270 67.700 ;
        RECT 14.430 67.250 17.260 67.300 ;
        RECT 14.310 67.130 17.260 67.250 ;
        RECT 14.310 65.720 14.600 67.130 ;
        RECT 14.940 66.260 15.110 66.590 ;
        RECT 15.325 66.560 16.365 66.730 ;
        RECT 15.325 66.120 16.365 66.290 ;
        RECT 16.580 66.260 16.750 66.590 ;
        RECT 17.090 65.720 17.260 67.130 ;
        RECT 14.310 65.600 17.260 65.720 ;
        RECT 14.430 65.550 17.260 65.600 ;
        RECT 17.820 67.220 20.560 67.290 ;
        RECT 21.140 67.220 23.880 67.290 ;
        RECT 17.820 67.120 20.690 67.220 ;
        RECT 17.820 65.710 17.990 67.120 ;
        RECT 18.330 66.250 18.500 66.580 ;
        RECT 18.670 66.550 19.710 66.720 ;
        RECT 18.670 66.110 19.710 66.280 ;
        RECT 19.880 66.250 20.050 66.580 ;
        RECT 20.390 65.710 20.690 67.120 ;
        RECT 17.820 65.570 20.690 65.710 ;
        RECT 21.010 67.120 23.880 67.220 ;
        RECT 21.010 65.710 21.310 67.120 ;
        RECT 21.650 66.250 21.820 66.580 ;
        RECT 21.990 66.550 23.030 66.720 ;
        RECT 21.990 66.110 23.030 66.280 ;
        RECT 23.200 66.250 23.370 66.580 ;
        RECT 23.710 65.710 23.880 67.120 ;
        RECT 21.010 65.570 23.880 65.710 ;
        RECT 17.820 65.540 20.560 65.570 ;
        RECT 21.140 65.540 23.880 65.570 ;
        RECT 24.440 67.250 27.270 67.300 ;
        RECT 24.440 67.130 27.390 67.250 ;
        RECT 24.440 65.720 24.610 67.130 ;
        RECT 24.950 66.260 25.120 66.590 ;
        RECT 25.335 66.560 26.375 66.730 ;
        RECT 25.335 66.120 26.375 66.290 ;
        RECT 26.590 66.260 26.760 66.590 ;
        RECT 27.100 65.720 27.390 67.130 ;
        RECT 24.440 65.600 27.390 65.720 ;
        RECT 24.440 65.550 27.270 65.600 ;
        RECT 14.430 65.150 17.260 65.200 ;
        RECT 14.310 65.030 17.260 65.150 ;
        RECT 14.310 63.620 14.600 65.030 ;
        RECT 14.940 64.160 15.110 64.490 ;
        RECT 15.325 64.460 16.365 64.630 ;
        RECT 15.325 64.020 16.365 64.190 ;
        RECT 16.580 64.160 16.750 64.490 ;
        RECT 17.090 63.620 17.260 65.030 ;
        RECT 14.310 63.500 17.260 63.620 ;
        RECT 14.430 63.450 17.260 63.500 ;
        RECT 17.820 65.120 20.560 65.190 ;
        RECT 21.140 65.120 23.880 65.190 ;
        RECT 17.820 65.020 20.690 65.120 ;
        RECT 17.820 63.610 17.990 65.020 ;
        RECT 18.330 64.150 18.500 64.480 ;
        RECT 18.670 64.450 19.710 64.620 ;
        RECT 18.670 64.010 19.710 64.180 ;
        RECT 19.880 64.150 20.050 64.480 ;
        RECT 20.390 63.610 20.690 65.020 ;
        RECT 17.820 63.470 20.690 63.610 ;
        RECT 21.010 65.020 23.880 65.120 ;
        RECT 21.010 63.610 21.310 65.020 ;
        RECT 21.650 64.150 21.820 64.480 ;
        RECT 21.990 64.450 23.030 64.620 ;
        RECT 21.990 64.010 23.030 64.180 ;
        RECT 23.200 64.150 23.370 64.480 ;
        RECT 23.710 63.610 23.880 65.020 ;
        RECT 21.010 63.470 23.880 63.610 ;
        RECT 17.820 63.440 20.560 63.470 ;
        RECT 21.140 63.440 23.880 63.470 ;
        RECT 24.440 65.150 27.270 65.200 ;
        RECT 24.440 65.030 27.390 65.150 ;
        RECT 24.440 63.620 24.610 65.030 ;
        RECT 24.950 64.160 25.120 64.490 ;
        RECT 25.335 64.460 26.375 64.630 ;
        RECT 25.335 64.020 26.375 64.190 ;
        RECT 26.590 64.160 26.760 64.490 ;
        RECT 27.100 63.620 27.390 65.030 ;
        RECT 24.440 63.500 27.390 63.620 ;
        RECT 24.440 63.450 27.270 63.500 ;
        RECT 14.430 63.050 17.260 63.100 ;
        RECT 14.310 62.930 17.260 63.050 ;
        RECT 14.310 61.520 14.600 62.930 ;
        RECT 14.940 62.060 15.110 62.390 ;
        RECT 15.325 62.360 16.365 62.530 ;
        RECT 15.325 61.920 16.365 62.090 ;
        RECT 16.580 62.060 16.750 62.390 ;
        RECT 17.090 61.520 17.260 62.930 ;
        RECT 14.310 61.400 17.260 61.520 ;
        RECT 14.430 61.350 17.260 61.400 ;
        RECT 17.820 63.020 20.560 63.090 ;
        RECT 21.140 63.020 23.880 63.090 ;
        RECT 17.820 62.920 20.690 63.020 ;
        RECT 17.820 61.510 17.990 62.920 ;
        RECT 18.330 62.050 18.500 62.380 ;
        RECT 18.670 62.350 19.710 62.520 ;
        RECT 18.670 61.910 19.710 62.080 ;
        RECT 19.880 62.050 20.050 62.380 ;
        RECT 20.390 61.510 20.690 62.920 ;
        RECT 17.820 61.370 20.690 61.510 ;
        RECT 21.010 62.920 23.880 63.020 ;
        RECT 21.010 61.510 21.310 62.920 ;
        RECT 21.650 62.050 21.820 62.380 ;
        RECT 21.990 62.350 23.030 62.520 ;
        RECT 21.990 61.910 23.030 62.080 ;
        RECT 23.200 62.050 23.370 62.380 ;
        RECT 23.710 61.510 23.880 62.920 ;
        RECT 21.010 61.370 23.880 61.510 ;
        RECT 17.820 61.340 20.560 61.370 ;
        RECT 21.140 61.340 23.880 61.370 ;
        RECT 24.440 63.050 27.270 63.100 ;
        RECT 24.440 62.930 27.390 63.050 ;
        RECT 24.440 61.520 24.610 62.930 ;
        RECT 24.950 62.060 25.120 62.390 ;
        RECT 25.335 62.360 26.375 62.530 ;
        RECT 25.335 61.920 26.375 62.090 ;
        RECT 26.590 62.060 26.760 62.390 ;
        RECT 27.100 61.520 27.390 62.930 ;
        RECT 24.440 61.400 27.390 61.520 ;
        RECT 24.440 61.350 27.270 61.400 ;
        RECT 14.430 60.950 17.260 61.000 ;
        RECT 14.310 60.830 17.260 60.950 ;
        RECT 14.310 59.420 14.600 60.830 ;
        RECT 14.940 59.960 15.110 60.290 ;
        RECT 15.325 60.260 16.365 60.430 ;
        RECT 15.325 59.820 16.365 59.990 ;
        RECT 16.580 59.960 16.750 60.290 ;
        RECT 17.090 59.420 17.260 60.830 ;
        RECT 14.310 59.300 17.260 59.420 ;
        RECT 14.430 59.250 17.260 59.300 ;
        RECT 17.820 60.920 20.560 60.990 ;
        RECT 21.140 60.920 23.880 60.990 ;
        RECT 17.820 60.820 20.690 60.920 ;
        RECT 17.820 59.410 17.990 60.820 ;
        RECT 18.330 59.950 18.500 60.280 ;
        RECT 18.670 60.250 19.710 60.420 ;
        RECT 18.670 59.810 19.710 59.980 ;
        RECT 19.880 59.950 20.050 60.280 ;
        RECT 20.390 59.410 20.690 60.820 ;
        RECT 17.820 59.270 20.690 59.410 ;
        RECT 21.010 60.820 23.880 60.920 ;
        RECT 21.010 59.410 21.310 60.820 ;
        RECT 21.650 59.950 21.820 60.280 ;
        RECT 21.990 60.250 23.030 60.420 ;
        RECT 21.990 59.810 23.030 59.980 ;
        RECT 23.200 59.950 23.370 60.280 ;
        RECT 23.710 59.410 23.880 60.820 ;
        RECT 21.010 59.270 23.880 59.410 ;
        RECT 17.820 59.240 20.560 59.270 ;
        RECT 21.140 59.240 23.880 59.270 ;
        RECT 24.440 60.950 27.270 61.000 ;
        RECT 24.440 60.830 27.390 60.950 ;
        RECT 24.440 59.420 24.610 60.830 ;
        RECT 24.950 59.960 25.120 60.290 ;
        RECT 25.335 60.260 26.375 60.430 ;
        RECT 25.335 59.820 26.375 59.990 ;
        RECT 26.590 59.960 26.760 60.290 ;
        RECT 27.100 59.420 27.390 60.830 ;
        RECT 24.440 59.300 27.390 59.420 ;
        RECT 24.440 59.250 27.270 59.300 ;
        RECT 14.430 58.850 17.260 58.900 ;
        RECT 14.310 58.730 17.260 58.850 ;
        RECT 14.310 57.320 14.600 58.730 ;
        RECT 14.940 57.860 15.110 58.190 ;
        RECT 15.325 58.160 16.365 58.330 ;
        RECT 15.325 57.720 16.365 57.890 ;
        RECT 16.580 57.860 16.750 58.190 ;
        RECT 17.090 57.320 17.260 58.730 ;
        RECT 14.310 57.200 17.260 57.320 ;
        RECT 14.430 57.150 17.260 57.200 ;
        RECT 17.820 58.820 20.560 58.890 ;
        RECT 21.140 58.820 23.880 58.890 ;
        RECT 17.820 58.720 20.690 58.820 ;
        RECT 17.820 57.310 17.990 58.720 ;
        RECT 18.330 57.850 18.500 58.180 ;
        RECT 18.670 58.150 19.710 58.320 ;
        RECT 18.670 57.710 19.710 57.880 ;
        RECT 19.880 57.850 20.050 58.180 ;
        RECT 20.390 57.310 20.690 58.720 ;
        RECT 17.820 57.170 20.690 57.310 ;
        RECT 21.010 58.720 23.880 58.820 ;
        RECT 21.010 57.310 21.310 58.720 ;
        RECT 21.650 57.850 21.820 58.180 ;
        RECT 21.990 58.150 23.030 58.320 ;
        RECT 21.990 57.710 23.030 57.880 ;
        RECT 23.200 57.850 23.370 58.180 ;
        RECT 23.710 57.310 23.880 58.720 ;
        RECT 21.010 57.170 23.880 57.310 ;
        RECT 17.820 57.140 20.560 57.170 ;
        RECT 21.140 57.140 23.880 57.170 ;
        RECT 24.440 58.850 27.270 58.900 ;
        RECT 24.440 58.730 27.390 58.850 ;
        RECT 24.440 57.320 24.610 58.730 ;
        RECT 24.950 57.860 25.120 58.190 ;
        RECT 25.335 58.160 26.375 58.330 ;
        RECT 25.335 57.720 26.375 57.890 ;
        RECT 26.590 57.860 26.760 58.190 ;
        RECT 27.100 57.320 27.390 58.730 ;
        RECT 24.440 57.200 27.390 57.320 ;
        RECT 24.440 57.150 27.270 57.200 ;
        RECT 14.430 56.750 17.260 56.800 ;
        RECT 14.310 56.630 17.260 56.750 ;
        RECT 14.310 55.220 14.600 56.630 ;
        RECT 14.940 55.760 15.110 56.090 ;
        RECT 15.325 56.060 16.365 56.230 ;
        RECT 15.325 55.620 16.365 55.790 ;
        RECT 16.580 55.760 16.750 56.090 ;
        RECT 17.090 55.220 17.260 56.630 ;
        RECT 14.310 55.100 17.260 55.220 ;
        RECT 14.430 55.050 17.260 55.100 ;
        RECT 17.820 56.720 20.560 56.790 ;
        RECT 21.140 56.720 23.880 56.790 ;
        RECT 17.820 56.620 20.690 56.720 ;
        RECT 17.820 55.210 17.990 56.620 ;
        RECT 18.330 55.750 18.500 56.080 ;
        RECT 18.670 56.050 19.710 56.220 ;
        RECT 18.670 55.610 19.710 55.780 ;
        RECT 19.880 55.750 20.050 56.080 ;
        RECT 20.390 55.210 20.690 56.620 ;
        RECT 17.820 55.070 20.690 55.210 ;
        RECT 21.010 56.620 23.880 56.720 ;
        RECT 21.010 55.210 21.310 56.620 ;
        RECT 21.650 55.750 21.820 56.080 ;
        RECT 21.990 56.050 23.030 56.220 ;
        RECT 21.990 55.610 23.030 55.780 ;
        RECT 23.200 55.750 23.370 56.080 ;
        RECT 23.710 55.210 23.880 56.620 ;
        RECT 21.010 55.070 23.880 55.210 ;
        RECT 17.820 55.040 20.560 55.070 ;
        RECT 21.140 55.040 23.880 55.070 ;
        RECT 24.440 56.750 27.270 56.800 ;
        RECT 24.440 56.630 27.390 56.750 ;
        RECT 24.440 55.220 24.610 56.630 ;
        RECT 24.950 55.760 25.120 56.090 ;
        RECT 25.335 56.060 26.375 56.230 ;
        RECT 25.335 55.620 26.375 55.790 ;
        RECT 26.590 55.760 26.760 56.090 ;
        RECT 27.100 55.220 27.390 56.630 ;
        RECT 24.440 55.100 27.390 55.220 ;
        RECT 24.440 55.050 27.270 55.100 ;
        RECT 14.430 54.650 17.260 54.700 ;
        RECT 14.310 54.530 17.260 54.650 ;
        RECT 14.310 53.120 14.600 54.530 ;
        RECT 14.940 53.660 15.110 53.990 ;
        RECT 15.325 53.960 16.365 54.130 ;
        RECT 15.325 53.520 16.365 53.690 ;
        RECT 16.580 53.660 16.750 53.990 ;
        RECT 17.090 53.120 17.260 54.530 ;
        RECT 14.310 53.000 17.260 53.120 ;
        RECT 14.430 52.950 17.260 53.000 ;
        RECT 17.820 54.620 20.560 54.690 ;
        RECT 21.140 54.620 23.880 54.690 ;
        RECT 17.820 54.520 20.690 54.620 ;
        RECT 17.820 53.110 17.990 54.520 ;
        RECT 18.330 53.650 18.500 53.980 ;
        RECT 18.670 53.950 19.710 54.120 ;
        RECT 18.670 53.510 19.710 53.680 ;
        RECT 19.880 53.650 20.050 53.980 ;
        RECT 20.390 53.110 20.690 54.520 ;
        RECT 17.820 52.970 20.690 53.110 ;
        RECT 21.010 54.520 23.880 54.620 ;
        RECT 21.010 53.110 21.310 54.520 ;
        RECT 21.650 53.650 21.820 53.980 ;
        RECT 21.990 53.950 23.030 54.120 ;
        RECT 21.990 53.510 23.030 53.680 ;
        RECT 23.200 53.650 23.370 53.980 ;
        RECT 23.710 53.110 23.880 54.520 ;
        RECT 21.010 52.970 23.880 53.110 ;
        RECT 17.820 52.940 20.560 52.970 ;
        RECT 21.140 52.940 23.880 52.970 ;
        RECT 24.440 54.650 27.270 54.700 ;
        RECT 24.440 54.530 27.390 54.650 ;
        RECT 24.440 53.120 24.610 54.530 ;
        RECT 24.950 53.660 25.120 53.990 ;
        RECT 25.335 53.960 26.375 54.130 ;
        RECT 25.335 53.520 26.375 53.690 ;
        RECT 26.590 53.660 26.760 53.990 ;
        RECT 27.100 53.120 27.390 54.530 ;
        RECT 24.440 53.000 27.390 53.120 ;
        RECT 24.440 52.950 27.270 53.000 ;
        RECT 14.430 52.550 17.260 52.600 ;
        RECT 14.310 52.430 17.260 52.550 ;
        RECT 14.310 51.020 14.600 52.430 ;
        RECT 14.940 51.560 15.110 51.890 ;
        RECT 15.325 51.860 16.365 52.030 ;
        RECT 15.325 51.420 16.365 51.590 ;
        RECT 16.580 51.560 16.750 51.890 ;
        RECT 17.090 51.020 17.260 52.430 ;
        RECT 14.310 50.900 17.260 51.020 ;
        RECT 14.430 50.850 17.260 50.900 ;
        RECT 17.820 52.520 20.560 52.590 ;
        RECT 21.140 52.520 23.880 52.590 ;
        RECT 17.820 52.420 20.690 52.520 ;
        RECT 17.820 51.010 17.990 52.420 ;
        RECT 18.330 51.550 18.500 51.880 ;
        RECT 18.670 51.850 19.710 52.020 ;
        RECT 18.670 51.410 19.710 51.580 ;
        RECT 19.880 51.550 20.050 51.880 ;
        RECT 20.390 51.010 20.690 52.420 ;
        RECT 17.820 50.870 20.690 51.010 ;
        RECT 21.010 52.420 23.880 52.520 ;
        RECT 21.010 51.010 21.310 52.420 ;
        RECT 21.650 51.550 21.820 51.880 ;
        RECT 21.990 51.850 23.030 52.020 ;
        RECT 21.990 51.410 23.030 51.580 ;
        RECT 23.200 51.550 23.370 51.880 ;
        RECT 23.710 51.010 23.880 52.420 ;
        RECT 21.010 50.870 23.880 51.010 ;
        RECT 17.820 50.840 20.560 50.870 ;
        RECT 21.140 50.840 23.880 50.870 ;
        RECT 24.440 52.550 27.270 52.600 ;
        RECT 24.440 52.430 27.390 52.550 ;
        RECT 24.440 51.020 24.610 52.430 ;
        RECT 24.950 51.560 25.120 51.890 ;
        RECT 25.335 51.860 26.375 52.030 ;
        RECT 25.335 51.420 26.375 51.590 ;
        RECT 26.590 51.560 26.760 51.890 ;
        RECT 27.100 51.020 27.390 52.430 ;
        RECT 24.440 50.900 27.390 51.020 ;
        RECT 24.440 50.850 27.270 50.900 ;
        RECT 14.430 50.450 17.260 50.500 ;
        RECT 14.310 50.330 17.260 50.450 ;
        RECT 14.310 48.920 14.600 50.330 ;
        RECT 14.940 49.460 15.110 49.790 ;
        RECT 15.325 49.760 16.365 49.930 ;
        RECT 15.325 49.320 16.365 49.490 ;
        RECT 16.580 49.460 16.750 49.790 ;
        RECT 17.090 48.920 17.260 50.330 ;
        RECT 14.310 48.800 17.260 48.920 ;
        RECT 14.430 48.750 17.260 48.800 ;
        RECT 17.820 50.420 20.560 50.490 ;
        RECT 21.140 50.420 23.880 50.490 ;
        RECT 17.820 50.320 20.690 50.420 ;
        RECT 17.820 48.910 17.990 50.320 ;
        RECT 18.330 49.450 18.500 49.780 ;
        RECT 18.670 49.750 19.710 49.920 ;
        RECT 18.670 49.310 19.710 49.480 ;
        RECT 19.880 49.450 20.050 49.780 ;
        RECT 20.390 48.910 20.690 50.320 ;
        RECT 17.820 48.770 20.690 48.910 ;
        RECT 21.010 50.320 23.880 50.420 ;
        RECT 21.010 48.910 21.310 50.320 ;
        RECT 21.650 49.450 21.820 49.780 ;
        RECT 21.990 49.750 23.030 49.920 ;
        RECT 21.990 49.310 23.030 49.480 ;
        RECT 23.200 49.450 23.370 49.780 ;
        RECT 23.710 48.910 23.880 50.320 ;
        RECT 21.010 48.770 23.880 48.910 ;
        RECT 17.820 48.740 20.560 48.770 ;
        RECT 21.140 48.740 23.880 48.770 ;
        RECT 24.440 50.450 27.270 50.500 ;
        RECT 24.440 50.330 27.390 50.450 ;
        RECT 24.440 48.920 24.610 50.330 ;
        RECT 24.950 49.460 25.120 49.790 ;
        RECT 25.335 49.760 26.375 49.930 ;
        RECT 25.335 49.320 26.375 49.490 ;
        RECT 26.590 49.460 26.760 49.790 ;
        RECT 27.100 48.920 27.390 50.330 ;
        RECT 24.440 48.800 27.390 48.920 ;
        RECT 24.440 48.750 27.270 48.800 ;
        RECT 14.430 48.350 17.260 48.400 ;
        RECT 14.310 48.230 17.260 48.350 ;
        RECT 14.310 46.820 14.600 48.230 ;
        RECT 14.940 47.360 15.110 47.690 ;
        RECT 15.325 47.660 16.365 47.830 ;
        RECT 15.325 47.220 16.365 47.390 ;
        RECT 16.580 47.360 16.750 47.690 ;
        RECT 17.090 46.820 17.260 48.230 ;
        RECT 14.310 46.700 17.260 46.820 ;
        RECT 14.430 46.650 17.260 46.700 ;
        RECT 17.820 48.320 20.560 48.390 ;
        RECT 21.140 48.320 23.880 48.390 ;
        RECT 17.820 48.220 20.690 48.320 ;
        RECT 17.820 46.810 17.990 48.220 ;
        RECT 18.330 47.350 18.500 47.680 ;
        RECT 18.670 47.650 19.710 47.820 ;
        RECT 18.670 47.210 19.710 47.380 ;
        RECT 19.880 47.350 20.050 47.680 ;
        RECT 20.390 46.810 20.690 48.220 ;
        RECT 17.820 46.670 20.690 46.810 ;
        RECT 21.010 48.220 23.880 48.320 ;
        RECT 21.010 46.810 21.310 48.220 ;
        RECT 21.650 47.350 21.820 47.680 ;
        RECT 21.990 47.650 23.030 47.820 ;
        RECT 21.990 47.210 23.030 47.380 ;
        RECT 23.200 47.350 23.370 47.680 ;
        RECT 23.710 46.810 23.880 48.220 ;
        RECT 21.010 46.670 23.880 46.810 ;
        RECT 17.820 46.640 20.560 46.670 ;
        RECT 21.140 46.640 23.880 46.670 ;
        RECT 24.440 48.350 27.270 48.400 ;
        RECT 24.440 48.230 27.390 48.350 ;
        RECT 24.440 46.820 24.610 48.230 ;
        RECT 24.950 47.360 25.120 47.690 ;
        RECT 25.335 47.660 26.375 47.830 ;
        RECT 25.335 47.220 26.375 47.390 ;
        RECT 26.590 47.360 26.760 47.690 ;
        RECT 27.100 46.820 27.390 48.230 ;
        RECT 24.440 46.700 27.390 46.820 ;
        RECT 24.440 46.650 27.270 46.700 ;
        RECT 14.430 46.250 17.260 46.300 ;
        RECT 14.310 46.130 17.260 46.250 ;
        RECT 14.310 44.720 14.600 46.130 ;
        RECT 14.940 45.260 15.110 45.590 ;
        RECT 15.325 45.560 16.365 45.730 ;
        RECT 15.325 45.120 16.365 45.290 ;
        RECT 16.580 45.260 16.750 45.590 ;
        RECT 17.090 44.720 17.260 46.130 ;
        RECT 14.310 44.600 17.260 44.720 ;
        RECT 14.430 44.550 17.260 44.600 ;
        RECT 17.820 46.220 20.560 46.290 ;
        RECT 21.140 46.220 23.880 46.290 ;
        RECT 17.820 46.120 20.690 46.220 ;
        RECT 17.820 44.710 17.990 46.120 ;
        RECT 18.330 45.250 18.500 45.580 ;
        RECT 18.670 45.550 19.710 45.720 ;
        RECT 18.670 45.110 19.710 45.280 ;
        RECT 19.880 45.250 20.050 45.580 ;
        RECT 20.390 44.710 20.690 46.120 ;
        RECT 17.820 44.570 20.690 44.710 ;
        RECT 21.010 46.120 23.880 46.220 ;
        RECT 21.010 44.710 21.310 46.120 ;
        RECT 21.650 45.250 21.820 45.580 ;
        RECT 21.990 45.550 23.030 45.720 ;
        RECT 21.990 45.110 23.030 45.280 ;
        RECT 23.200 45.250 23.370 45.580 ;
        RECT 23.710 44.710 23.880 46.120 ;
        RECT 21.010 44.570 23.880 44.710 ;
        RECT 17.820 44.540 20.560 44.570 ;
        RECT 21.140 44.540 23.880 44.570 ;
        RECT 24.440 46.250 27.270 46.300 ;
        RECT 24.440 46.130 27.390 46.250 ;
        RECT 24.440 44.720 24.610 46.130 ;
        RECT 24.950 45.260 25.120 45.590 ;
        RECT 25.335 45.560 26.375 45.730 ;
        RECT 25.335 45.120 26.375 45.290 ;
        RECT 26.590 45.260 26.760 45.590 ;
        RECT 27.100 44.720 27.390 46.130 ;
        RECT 24.440 44.600 27.390 44.720 ;
        RECT 24.440 44.550 27.270 44.600 ;
        RECT 14.430 44.150 17.260 44.200 ;
        RECT 14.310 44.030 17.260 44.150 ;
        RECT 14.310 42.620 14.600 44.030 ;
        RECT 14.940 43.160 15.110 43.490 ;
        RECT 15.325 43.460 16.365 43.630 ;
        RECT 15.325 43.020 16.365 43.190 ;
        RECT 16.580 43.160 16.750 43.490 ;
        RECT 17.090 42.620 17.260 44.030 ;
        RECT 14.310 42.500 17.260 42.620 ;
        RECT 14.430 42.450 17.260 42.500 ;
        RECT 17.820 44.120 20.560 44.190 ;
        RECT 21.140 44.120 23.880 44.190 ;
        RECT 17.820 44.020 20.690 44.120 ;
        RECT 17.820 42.610 17.990 44.020 ;
        RECT 18.330 43.150 18.500 43.480 ;
        RECT 18.670 43.450 19.710 43.620 ;
        RECT 18.670 43.010 19.710 43.180 ;
        RECT 19.880 43.150 20.050 43.480 ;
        RECT 20.390 42.610 20.690 44.020 ;
        RECT 17.820 42.470 20.690 42.610 ;
        RECT 21.010 44.020 23.880 44.120 ;
        RECT 21.010 42.610 21.310 44.020 ;
        RECT 21.650 43.150 21.820 43.480 ;
        RECT 21.990 43.450 23.030 43.620 ;
        RECT 21.990 43.010 23.030 43.180 ;
        RECT 23.200 43.150 23.370 43.480 ;
        RECT 23.710 42.610 23.880 44.020 ;
        RECT 21.010 42.470 23.880 42.610 ;
        RECT 17.820 42.440 20.560 42.470 ;
        RECT 21.140 42.440 23.880 42.470 ;
        RECT 24.440 44.150 27.270 44.200 ;
        RECT 24.440 44.030 27.390 44.150 ;
        RECT 24.440 42.620 24.610 44.030 ;
        RECT 24.950 43.160 25.120 43.490 ;
        RECT 25.335 43.460 26.375 43.630 ;
        RECT 25.335 43.020 26.375 43.190 ;
        RECT 26.590 43.160 26.760 43.490 ;
        RECT 27.100 42.620 27.390 44.030 ;
        RECT 24.440 42.500 27.390 42.620 ;
        RECT 24.440 42.450 27.270 42.500 ;
        RECT 14.430 42.050 17.260 42.100 ;
        RECT 14.310 41.930 17.260 42.050 ;
        RECT 14.310 40.520 14.600 41.930 ;
        RECT 14.940 41.060 15.110 41.390 ;
        RECT 15.325 41.360 16.365 41.530 ;
        RECT 15.325 40.920 16.365 41.090 ;
        RECT 16.580 41.060 16.750 41.390 ;
        RECT 17.090 40.520 17.260 41.930 ;
        RECT 14.310 40.400 17.260 40.520 ;
        RECT 14.430 40.350 17.260 40.400 ;
        RECT 17.820 42.020 20.560 42.090 ;
        RECT 21.140 42.020 23.880 42.090 ;
        RECT 17.820 41.920 20.690 42.020 ;
        RECT 17.820 40.510 17.990 41.920 ;
        RECT 18.330 41.050 18.500 41.380 ;
        RECT 18.670 41.350 19.710 41.520 ;
        RECT 18.670 40.910 19.710 41.080 ;
        RECT 19.880 41.050 20.050 41.380 ;
        RECT 20.390 40.510 20.690 41.920 ;
        RECT 17.820 40.370 20.690 40.510 ;
        RECT 21.010 41.920 23.880 42.020 ;
        RECT 21.010 40.510 21.310 41.920 ;
        RECT 21.650 41.050 21.820 41.380 ;
        RECT 21.990 41.350 23.030 41.520 ;
        RECT 21.990 40.910 23.030 41.080 ;
        RECT 23.200 41.050 23.370 41.380 ;
        RECT 23.710 40.510 23.880 41.920 ;
        RECT 21.010 40.370 23.880 40.510 ;
        RECT 17.820 40.340 20.560 40.370 ;
        RECT 21.140 40.340 23.880 40.370 ;
        RECT 24.440 42.050 27.270 42.100 ;
        RECT 24.440 41.930 27.390 42.050 ;
        RECT 24.440 40.520 24.610 41.930 ;
        RECT 24.950 41.060 25.120 41.390 ;
        RECT 25.335 41.360 26.375 41.530 ;
        RECT 25.335 40.920 26.375 41.090 ;
        RECT 26.590 41.060 26.760 41.390 ;
        RECT 27.100 40.520 27.390 41.930 ;
        RECT 24.440 40.400 27.390 40.520 ;
        RECT 24.440 40.350 27.270 40.400 ;
        RECT 14.430 39.950 17.260 40.000 ;
        RECT 14.310 39.830 17.260 39.950 ;
        RECT 14.310 38.420 14.600 39.830 ;
        RECT 14.940 38.960 15.110 39.290 ;
        RECT 15.325 39.260 16.365 39.430 ;
        RECT 15.325 38.820 16.365 38.990 ;
        RECT 16.580 38.960 16.750 39.290 ;
        RECT 17.090 38.420 17.260 39.830 ;
        RECT 14.310 38.300 17.260 38.420 ;
        RECT 14.430 38.250 17.260 38.300 ;
        RECT 17.820 39.920 20.560 39.990 ;
        RECT 21.140 39.920 23.880 39.990 ;
        RECT 17.820 39.820 20.690 39.920 ;
        RECT 17.820 38.410 17.990 39.820 ;
        RECT 18.330 38.950 18.500 39.280 ;
        RECT 18.670 39.250 19.710 39.420 ;
        RECT 18.670 38.810 19.710 38.980 ;
        RECT 19.880 38.950 20.050 39.280 ;
        RECT 20.390 38.410 20.690 39.820 ;
        RECT 17.820 38.270 20.690 38.410 ;
        RECT 21.010 39.820 23.880 39.920 ;
        RECT 21.010 38.410 21.310 39.820 ;
        RECT 21.650 38.950 21.820 39.280 ;
        RECT 21.990 39.250 23.030 39.420 ;
        RECT 21.990 38.810 23.030 38.980 ;
        RECT 23.200 38.950 23.370 39.280 ;
        RECT 23.710 38.410 23.880 39.820 ;
        RECT 21.010 38.270 23.880 38.410 ;
        RECT 17.820 38.240 20.560 38.270 ;
        RECT 21.140 38.240 23.880 38.270 ;
        RECT 24.440 39.950 27.270 40.000 ;
        RECT 24.440 39.830 27.390 39.950 ;
        RECT 24.440 38.420 24.610 39.830 ;
        RECT 24.950 38.960 25.120 39.290 ;
        RECT 25.335 39.260 26.375 39.430 ;
        RECT 25.335 38.820 26.375 38.990 ;
        RECT 26.590 38.960 26.760 39.290 ;
        RECT 27.100 38.420 27.390 39.830 ;
        RECT 24.440 38.300 27.390 38.420 ;
        RECT 24.440 38.250 27.270 38.300 ;
        RECT 14.430 37.850 17.260 37.900 ;
        RECT 14.310 37.730 17.260 37.850 ;
        RECT 14.310 36.320 14.600 37.730 ;
        RECT 14.940 36.860 15.110 37.190 ;
        RECT 15.325 37.160 16.365 37.330 ;
        RECT 15.325 36.720 16.365 36.890 ;
        RECT 16.580 36.860 16.750 37.190 ;
        RECT 17.090 36.320 17.260 37.730 ;
        RECT 14.310 36.200 17.260 36.320 ;
        RECT 14.430 36.150 17.260 36.200 ;
        RECT 17.820 37.820 20.560 37.890 ;
        RECT 21.140 37.820 23.880 37.890 ;
        RECT 17.820 37.720 20.690 37.820 ;
        RECT 17.820 36.310 17.990 37.720 ;
        RECT 18.330 36.850 18.500 37.180 ;
        RECT 18.670 37.150 19.710 37.320 ;
        RECT 18.670 36.710 19.710 36.880 ;
        RECT 19.880 36.850 20.050 37.180 ;
        RECT 20.390 36.310 20.690 37.720 ;
        RECT 17.820 36.170 20.690 36.310 ;
        RECT 21.010 37.720 23.880 37.820 ;
        RECT 21.010 36.310 21.310 37.720 ;
        RECT 21.650 36.850 21.820 37.180 ;
        RECT 21.990 37.150 23.030 37.320 ;
        RECT 21.990 36.710 23.030 36.880 ;
        RECT 23.200 36.850 23.370 37.180 ;
        RECT 23.710 36.310 23.880 37.720 ;
        RECT 21.010 36.170 23.880 36.310 ;
        RECT 17.820 36.140 20.560 36.170 ;
        RECT 21.140 36.140 23.880 36.170 ;
        RECT 24.440 37.850 27.270 37.900 ;
        RECT 24.440 37.730 27.390 37.850 ;
        RECT 24.440 36.320 24.610 37.730 ;
        RECT 24.950 36.860 25.120 37.190 ;
        RECT 25.335 37.160 26.375 37.330 ;
        RECT 25.335 36.720 26.375 36.890 ;
        RECT 26.590 36.860 26.760 37.190 ;
        RECT 27.100 36.320 27.390 37.730 ;
        RECT 24.440 36.200 27.390 36.320 ;
        RECT 24.440 36.150 27.270 36.200 ;
        RECT 14.430 35.750 17.260 35.800 ;
        RECT 14.310 35.630 17.260 35.750 ;
        RECT 14.310 34.220 14.600 35.630 ;
        RECT 14.940 34.760 15.110 35.090 ;
        RECT 15.325 35.060 16.365 35.230 ;
        RECT 15.325 34.620 16.365 34.790 ;
        RECT 16.580 34.760 16.750 35.090 ;
        RECT 17.090 34.220 17.260 35.630 ;
        RECT 14.310 34.100 17.260 34.220 ;
        RECT 14.430 34.050 17.260 34.100 ;
        RECT 17.820 35.720 20.560 35.790 ;
        RECT 21.140 35.720 23.880 35.790 ;
        RECT 17.820 35.620 20.690 35.720 ;
        RECT 17.820 34.210 17.990 35.620 ;
        RECT 18.330 34.750 18.500 35.080 ;
        RECT 18.670 35.050 19.710 35.220 ;
        RECT 18.670 34.610 19.710 34.780 ;
        RECT 19.880 34.750 20.050 35.080 ;
        RECT 20.390 34.210 20.690 35.620 ;
        RECT 17.820 34.070 20.690 34.210 ;
        RECT 21.010 35.620 23.880 35.720 ;
        RECT 21.010 34.210 21.310 35.620 ;
        RECT 21.650 34.750 21.820 35.080 ;
        RECT 21.990 35.050 23.030 35.220 ;
        RECT 21.990 34.610 23.030 34.780 ;
        RECT 23.200 34.750 23.370 35.080 ;
        RECT 23.710 34.210 23.880 35.620 ;
        RECT 21.010 34.070 23.880 34.210 ;
        RECT 17.820 34.040 20.560 34.070 ;
        RECT 21.140 34.040 23.880 34.070 ;
        RECT 24.440 35.750 27.270 35.800 ;
        RECT 24.440 35.630 27.390 35.750 ;
        RECT 24.440 34.220 24.610 35.630 ;
        RECT 24.950 34.760 25.120 35.090 ;
        RECT 25.335 35.060 26.375 35.230 ;
        RECT 25.335 34.620 26.375 34.790 ;
        RECT 26.590 34.760 26.760 35.090 ;
        RECT 27.100 34.220 27.390 35.630 ;
        RECT 24.440 34.100 27.390 34.220 ;
        RECT 24.440 34.050 27.270 34.100 ;
        RECT 14.430 33.650 17.260 33.700 ;
        RECT 14.310 33.530 17.260 33.650 ;
        RECT 14.310 32.120 14.600 33.530 ;
        RECT 14.940 32.660 15.110 32.990 ;
        RECT 15.325 32.960 16.365 33.130 ;
        RECT 15.325 32.520 16.365 32.690 ;
        RECT 16.580 32.660 16.750 32.990 ;
        RECT 17.090 32.120 17.260 33.530 ;
        RECT 14.310 32.000 17.260 32.120 ;
        RECT 14.430 31.950 17.260 32.000 ;
        RECT 17.820 33.620 20.560 33.690 ;
        RECT 21.140 33.620 23.880 33.690 ;
        RECT 17.820 33.520 20.690 33.620 ;
        RECT 17.820 32.110 17.990 33.520 ;
        RECT 18.330 32.650 18.500 32.980 ;
        RECT 18.670 32.950 19.710 33.120 ;
        RECT 18.670 32.510 19.710 32.680 ;
        RECT 19.880 32.650 20.050 32.980 ;
        RECT 20.390 32.110 20.690 33.520 ;
        RECT 17.820 31.970 20.690 32.110 ;
        RECT 21.010 33.520 23.880 33.620 ;
        RECT 21.010 32.110 21.310 33.520 ;
        RECT 21.650 32.650 21.820 32.980 ;
        RECT 21.990 32.950 23.030 33.120 ;
        RECT 21.990 32.510 23.030 32.680 ;
        RECT 23.200 32.650 23.370 32.980 ;
        RECT 23.710 32.110 23.880 33.520 ;
        RECT 21.010 31.970 23.880 32.110 ;
        RECT 17.820 31.940 20.560 31.970 ;
        RECT 21.140 31.940 23.880 31.970 ;
        RECT 24.440 33.650 27.270 33.700 ;
        RECT 24.440 33.530 27.390 33.650 ;
        RECT 24.440 32.120 24.610 33.530 ;
        RECT 24.950 32.660 25.120 32.990 ;
        RECT 25.335 32.960 26.375 33.130 ;
        RECT 25.335 32.520 26.375 32.690 ;
        RECT 26.590 32.660 26.760 32.990 ;
        RECT 27.100 32.120 27.390 33.530 ;
        RECT 24.440 32.000 27.390 32.120 ;
        RECT 24.440 31.950 27.270 32.000 ;
        RECT 14.430 31.550 17.260 31.600 ;
        RECT 14.310 31.430 17.260 31.550 ;
        RECT 14.310 30.020 14.600 31.430 ;
        RECT 14.940 30.560 15.110 30.890 ;
        RECT 15.325 30.860 16.365 31.030 ;
        RECT 15.325 30.420 16.365 30.590 ;
        RECT 16.580 30.560 16.750 30.890 ;
        RECT 17.090 30.020 17.260 31.430 ;
        RECT 14.310 29.900 17.260 30.020 ;
        RECT 14.430 29.850 17.260 29.900 ;
        RECT 17.820 31.520 20.560 31.590 ;
        RECT 21.140 31.520 23.880 31.590 ;
        RECT 17.820 31.420 20.690 31.520 ;
        RECT 17.820 30.010 17.990 31.420 ;
        RECT 18.330 30.550 18.500 30.880 ;
        RECT 18.670 30.850 19.710 31.020 ;
        RECT 18.670 30.410 19.710 30.580 ;
        RECT 19.880 30.550 20.050 30.880 ;
        RECT 20.390 30.010 20.690 31.420 ;
        RECT 17.820 29.870 20.690 30.010 ;
        RECT 21.010 31.420 23.880 31.520 ;
        RECT 21.010 30.010 21.310 31.420 ;
        RECT 21.650 30.550 21.820 30.880 ;
        RECT 21.990 30.850 23.030 31.020 ;
        RECT 21.990 30.410 23.030 30.580 ;
        RECT 23.200 30.550 23.370 30.880 ;
        RECT 23.710 30.010 23.880 31.420 ;
        RECT 21.010 29.870 23.880 30.010 ;
        RECT 17.820 29.840 20.560 29.870 ;
        RECT 21.140 29.840 23.880 29.870 ;
        RECT 24.440 31.550 27.270 31.600 ;
        RECT 24.440 31.430 27.390 31.550 ;
        RECT 24.440 30.020 24.610 31.430 ;
        RECT 24.950 30.560 25.120 30.890 ;
        RECT 25.335 30.860 26.375 31.030 ;
        RECT 25.335 30.420 26.375 30.590 ;
        RECT 26.590 30.560 26.760 30.890 ;
        RECT 27.100 30.020 27.390 31.430 ;
        RECT 24.440 29.900 27.390 30.020 ;
        RECT 24.440 29.850 27.270 29.900 ;
        RECT 14.430 29.450 17.260 29.500 ;
        RECT 14.310 29.330 17.260 29.450 ;
        RECT 14.310 27.920 14.600 29.330 ;
        RECT 14.940 28.460 15.110 28.790 ;
        RECT 15.325 28.760 16.365 28.930 ;
        RECT 15.325 28.320 16.365 28.490 ;
        RECT 16.580 28.460 16.750 28.790 ;
        RECT 17.090 27.920 17.260 29.330 ;
        RECT 14.310 27.800 17.260 27.920 ;
        RECT 14.430 27.750 17.260 27.800 ;
        RECT 17.820 29.420 20.560 29.490 ;
        RECT 21.140 29.420 23.880 29.490 ;
        RECT 17.820 29.320 20.690 29.420 ;
        RECT 17.820 27.910 17.990 29.320 ;
        RECT 18.330 28.450 18.500 28.780 ;
        RECT 18.670 28.750 19.710 28.920 ;
        RECT 18.670 28.310 19.710 28.480 ;
        RECT 19.880 28.450 20.050 28.780 ;
        RECT 20.390 27.910 20.690 29.320 ;
        RECT 17.820 27.770 20.690 27.910 ;
        RECT 21.010 29.320 23.880 29.420 ;
        RECT 21.010 27.910 21.310 29.320 ;
        RECT 21.650 28.450 21.820 28.780 ;
        RECT 21.990 28.750 23.030 28.920 ;
        RECT 21.990 28.310 23.030 28.480 ;
        RECT 23.200 28.450 23.370 28.780 ;
        RECT 23.710 27.910 23.880 29.320 ;
        RECT 21.010 27.770 23.880 27.910 ;
        RECT 17.820 27.740 20.560 27.770 ;
        RECT 21.140 27.740 23.880 27.770 ;
        RECT 24.440 29.450 27.270 29.500 ;
        RECT 24.440 29.330 27.390 29.450 ;
        RECT 24.440 27.920 24.610 29.330 ;
        RECT 24.950 28.460 25.120 28.790 ;
        RECT 25.335 28.760 26.375 28.930 ;
        RECT 25.335 28.320 26.375 28.490 ;
        RECT 26.590 28.460 26.760 28.790 ;
        RECT 27.100 27.920 27.390 29.330 ;
        RECT 24.440 27.800 27.390 27.920 ;
        RECT 24.440 27.750 27.270 27.800 ;
        RECT 14.430 27.350 17.260 27.400 ;
        RECT 14.310 27.230 17.260 27.350 ;
        RECT 14.310 25.820 14.600 27.230 ;
        RECT 14.940 26.360 15.110 26.690 ;
        RECT 15.325 26.660 16.365 26.830 ;
        RECT 15.325 26.220 16.365 26.390 ;
        RECT 16.580 26.360 16.750 26.690 ;
        RECT 17.090 25.820 17.260 27.230 ;
        RECT 14.310 25.700 17.260 25.820 ;
        RECT 14.430 25.650 17.260 25.700 ;
        RECT 17.820 27.320 20.560 27.390 ;
        RECT 21.140 27.320 23.880 27.390 ;
        RECT 17.820 27.220 20.690 27.320 ;
        RECT 17.820 25.810 17.990 27.220 ;
        RECT 18.330 26.350 18.500 26.680 ;
        RECT 18.670 26.650 19.710 26.820 ;
        RECT 18.670 26.210 19.710 26.380 ;
        RECT 19.880 26.350 20.050 26.680 ;
        RECT 20.390 25.810 20.690 27.220 ;
        RECT 17.820 25.670 20.690 25.810 ;
        RECT 21.010 27.220 23.880 27.320 ;
        RECT 21.010 25.810 21.310 27.220 ;
        RECT 21.650 26.350 21.820 26.680 ;
        RECT 21.990 26.650 23.030 26.820 ;
        RECT 21.990 26.210 23.030 26.380 ;
        RECT 23.200 26.350 23.370 26.680 ;
        RECT 23.710 25.810 23.880 27.220 ;
        RECT 21.010 25.670 23.880 25.810 ;
        RECT 17.820 25.640 20.560 25.670 ;
        RECT 21.140 25.640 23.880 25.670 ;
        RECT 24.440 27.350 27.270 27.400 ;
        RECT 24.440 27.230 27.390 27.350 ;
        RECT 24.440 25.820 24.610 27.230 ;
        RECT 24.950 26.360 25.120 26.690 ;
        RECT 25.335 26.660 26.375 26.830 ;
        RECT 25.335 26.220 26.375 26.390 ;
        RECT 26.590 26.360 26.760 26.690 ;
        RECT 27.100 25.820 27.390 27.230 ;
        RECT 24.440 25.700 27.390 25.820 ;
        RECT 24.440 25.650 27.270 25.700 ;
        RECT 14.430 25.250 17.260 25.300 ;
        RECT 14.310 25.130 17.260 25.250 ;
        RECT 14.310 23.720 14.600 25.130 ;
        RECT 14.940 24.260 15.110 24.590 ;
        RECT 15.325 24.560 16.365 24.730 ;
        RECT 15.325 24.120 16.365 24.290 ;
        RECT 16.580 24.260 16.750 24.590 ;
        RECT 17.090 23.720 17.260 25.130 ;
        RECT 14.310 23.600 17.260 23.720 ;
        RECT 14.430 23.550 17.260 23.600 ;
        RECT 17.820 25.220 20.560 25.290 ;
        RECT 21.140 25.220 23.880 25.290 ;
        RECT 17.820 25.120 20.690 25.220 ;
        RECT 17.820 23.710 17.990 25.120 ;
        RECT 18.330 24.250 18.500 24.580 ;
        RECT 18.670 24.550 19.710 24.720 ;
        RECT 18.670 24.110 19.710 24.280 ;
        RECT 19.880 24.250 20.050 24.580 ;
        RECT 20.390 23.710 20.690 25.120 ;
        RECT 17.820 23.570 20.690 23.710 ;
        RECT 21.010 25.120 23.880 25.220 ;
        RECT 21.010 23.710 21.310 25.120 ;
        RECT 21.650 24.250 21.820 24.580 ;
        RECT 21.990 24.550 23.030 24.720 ;
        RECT 21.990 24.110 23.030 24.280 ;
        RECT 23.200 24.250 23.370 24.580 ;
        RECT 23.710 23.710 23.880 25.120 ;
        RECT 21.010 23.570 23.880 23.710 ;
        RECT 17.820 23.540 20.560 23.570 ;
        RECT 21.140 23.540 23.880 23.570 ;
        RECT 24.440 25.250 27.270 25.300 ;
        RECT 24.440 25.130 27.390 25.250 ;
        RECT 24.440 23.720 24.610 25.130 ;
        RECT 24.950 24.260 25.120 24.590 ;
        RECT 25.335 24.560 26.375 24.730 ;
        RECT 25.335 24.120 26.375 24.290 ;
        RECT 26.590 24.260 26.760 24.590 ;
        RECT 27.100 23.720 27.390 25.130 ;
        RECT 24.440 23.600 27.390 23.720 ;
        RECT 24.440 23.550 27.270 23.600 ;
        RECT 14.430 23.150 17.260 23.200 ;
        RECT 14.310 23.030 17.260 23.150 ;
        RECT 14.310 21.620 14.600 23.030 ;
        RECT 14.940 22.160 15.110 22.490 ;
        RECT 15.325 22.460 16.365 22.630 ;
        RECT 15.325 22.020 16.365 22.190 ;
        RECT 16.580 22.160 16.750 22.490 ;
        RECT 17.090 21.620 17.260 23.030 ;
        RECT 14.310 21.500 17.260 21.620 ;
        RECT 14.430 21.450 17.260 21.500 ;
        RECT 17.820 23.120 20.560 23.190 ;
        RECT 21.140 23.120 23.880 23.190 ;
        RECT 17.820 23.020 20.690 23.120 ;
        RECT 17.820 21.610 17.990 23.020 ;
        RECT 18.330 22.150 18.500 22.480 ;
        RECT 18.670 22.450 19.710 22.620 ;
        RECT 18.670 22.010 19.710 22.180 ;
        RECT 19.880 22.150 20.050 22.480 ;
        RECT 20.390 21.610 20.690 23.020 ;
        RECT 17.820 21.470 20.690 21.610 ;
        RECT 21.010 23.020 23.880 23.120 ;
        RECT 21.010 21.610 21.310 23.020 ;
        RECT 21.650 22.150 21.820 22.480 ;
        RECT 21.990 22.450 23.030 22.620 ;
        RECT 21.990 22.010 23.030 22.180 ;
        RECT 23.200 22.150 23.370 22.480 ;
        RECT 23.710 21.610 23.880 23.020 ;
        RECT 21.010 21.470 23.880 21.610 ;
        RECT 17.820 21.440 20.560 21.470 ;
        RECT 21.140 21.440 23.880 21.470 ;
        RECT 24.440 23.150 27.270 23.200 ;
        RECT 24.440 23.030 27.390 23.150 ;
        RECT 24.440 21.620 24.610 23.030 ;
        RECT 24.950 22.160 25.120 22.490 ;
        RECT 25.335 22.460 26.375 22.630 ;
        RECT 25.335 22.020 26.375 22.190 ;
        RECT 26.590 22.160 26.760 22.490 ;
        RECT 27.100 21.620 27.390 23.030 ;
        RECT 24.440 21.500 27.390 21.620 ;
        RECT 24.440 21.450 27.270 21.500 ;
        RECT 14.430 21.050 17.260 21.100 ;
        RECT 14.310 20.930 17.260 21.050 ;
        RECT 14.310 19.520 14.600 20.930 ;
        RECT 14.940 20.060 15.110 20.390 ;
        RECT 15.325 20.360 16.365 20.530 ;
        RECT 15.325 19.920 16.365 20.090 ;
        RECT 16.580 20.060 16.750 20.390 ;
        RECT 17.090 19.520 17.260 20.930 ;
        RECT 14.310 19.400 17.260 19.520 ;
        RECT 14.430 19.350 17.260 19.400 ;
        RECT 17.820 21.020 20.560 21.090 ;
        RECT 21.140 21.020 23.880 21.090 ;
        RECT 17.820 20.920 20.690 21.020 ;
        RECT 17.820 19.510 17.990 20.920 ;
        RECT 18.330 20.050 18.500 20.380 ;
        RECT 18.670 20.350 19.710 20.520 ;
        RECT 18.670 19.910 19.710 20.080 ;
        RECT 19.880 20.050 20.050 20.380 ;
        RECT 20.390 19.510 20.690 20.920 ;
        RECT 17.820 19.370 20.690 19.510 ;
        RECT 21.010 20.920 23.880 21.020 ;
        RECT 21.010 19.510 21.310 20.920 ;
        RECT 21.650 20.050 21.820 20.380 ;
        RECT 21.990 20.350 23.030 20.520 ;
        RECT 21.990 19.910 23.030 20.080 ;
        RECT 23.200 20.050 23.370 20.380 ;
        RECT 23.710 19.510 23.880 20.920 ;
        RECT 21.010 19.370 23.880 19.510 ;
        RECT 17.820 19.340 20.560 19.370 ;
        RECT 21.140 19.340 23.880 19.370 ;
        RECT 24.440 21.050 27.270 21.100 ;
        RECT 24.440 20.930 27.390 21.050 ;
        RECT 24.440 19.520 24.610 20.930 ;
        RECT 24.950 20.060 25.120 20.390 ;
        RECT 25.335 20.360 26.375 20.530 ;
        RECT 25.335 19.920 26.375 20.090 ;
        RECT 26.590 20.060 26.760 20.390 ;
        RECT 27.100 19.520 27.390 20.930 ;
        RECT 24.440 19.400 27.390 19.520 ;
        RECT 24.440 19.350 27.270 19.400 ;
        RECT 14.430 18.950 17.260 19.000 ;
        RECT 14.310 18.830 17.260 18.950 ;
        RECT 14.310 17.420 14.600 18.830 ;
        RECT 14.940 17.960 15.110 18.290 ;
        RECT 15.325 18.260 16.365 18.430 ;
        RECT 15.325 17.820 16.365 17.990 ;
        RECT 16.580 17.960 16.750 18.290 ;
        RECT 17.090 17.420 17.260 18.830 ;
        RECT 14.310 17.300 17.260 17.420 ;
        RECT 14.430 17.250 17.260 17.300 ;
        RECT 17.820 18.920 20.560 18.990 ;
        RECT 21.140 18.920 23.880 18.990 ;
        RECT 17.820 18.820 20.690 18.920 ;
        RECT 17.820 17.410 17.990 18.820 ;
        RECT 18.330 17.950 18.500 18.280 ;
        RECT 18.670 18.250 19.710 18.420 ;
        RECT 18.670 17.810 19.710 17.980 ;
        RECT 19.880 17.950 20.050 18.280 ;
        RECT 20.390 17.410 20.690 18.820 ;
        RECT 17.820 17.270 20.690 17.410 ;
        RECT 21.010 18.820 23.880 18.920 ;
        RECT 21.010 17.410 21.310 18.820 ;
        RECT 21.650 17.950 21.820 18.280 ;
        RECT 21.990 18.250 23.030 18.420 ;
        RECT 21.990 17.810 23.030 17.980 ;
        RECT 23.200 17.950 23.370 18.280 ;
        RECT 23.710 17.410 23.880 18.820 ;
        RECT 21.010 17.270 23.880 17.410 ;
        RECT 17.820 17.240 20.560 17.270 ;
        RECT 21.140 17.240 23.880 17.270 ;
        RECT 24.440 18.950 27.270 19.000 ;
        RECT 24.440 18.830 27.390 18.950 ;
        RECT 24.440 17.420 24.610 18.830 ;
        RECT 24.950 17.960 25.120 18.290 ;
        RECT 25.335 18.260 26.375 18.430 ;
        RECT 25.335 17.820 26.375 17.990 ;
        RECT 26.590 17.960 26.760 18.290 ;
        RECT 27.100 17.420 27.390 18.830 ;
        RECT 24.440 17.300 27.390 17.420 ;
        RECT 24.440 17.250 27.270 17.300 ;
        RECT 14.430 16.850 17.260 16.900 ;
        RECT 14.310 16.730 17.260 16.850 ;
        RECT 14.310 15.320 14.600 16.730 ;
        RECT 14.940 15.860 15.110 16.190 ;
        RECT 15.325 16.160 16.365 16.330 ;
        RECT 15.325 15.720 16.365 15.890 ;
        RECT 16.580 15.860 16.750 16.190 ;
        RECT 17.090 15.320 17.260 16.730 ;
        RECT 14.310 15.200 17.260 15.320 ;
        RECT 14.430 15.150 17.260 15.200 ;
        RECT 17.820 16.820 20.560 16.890 ;
        RECT 21.140 16.820 23.880 16.890 ;
        RECT 17.820 16.720 20.690 16.820 ;
        RECT 17.820 15.310 17.990 16.720 ;
        RECT 18.330 15.850 18.500 16.180 ;
        RECT 18.670 16.150 19.710 16.320 ;
        RECT 18.670 15.710 19.710 15.880 ;
        RECT 19.880 15.850 20.050 16.180 ;
        RECT 20.390 15.310 20.690 16.720 ;
        RECT 17.820 15.170 20.690 15.310 ;
        RECT 21.010 16.720 23.880 16.820 ;
        RECT 21.010 15.310 21.310 16.720 ;
        RECT 21.650 15.850 21.820 16.180 ;
        RECT 21.990 16.150 23.030 16.320 ;
        RECT 21.990 15.710 23.030 15.880 ;
        RECT 23.200 15.850 23.370 16.180 ;
        RECT 23.710 15.310 23.880 16.720 ;
        RECT 21.010 15.170 23.880 15.310 ;
        RECT 17.820 15.140 20.560 15.170 ;
        RECT 21.140 15.140 23.880 15.170 ;
        RECT 24.440 16.850 27.270 16.900 ;
        RECT 24.440 16.730 27.390 16.850 ;
        RECT 24.440 15.320 24.610 16.730 ;
        RECT 24.950 15.860 25.120 16.190 ;
        RECT 25.335 16.160 26.375 16.330 ;
        RECT 25.335 15.720 26.375 15.890 ;
        RECT 26.590 15.860 26.760 16.190 ;
        RECT 27.100 15.320 27.390 16.730 ;
        RECT 24.440 15.200 27.390 15.320 ;
        RECT 24.440 15.150 27.270 15.200 ;
        RECT 14.430 14.750 17.260 14.800 ;
        RECT 14.310 14.630 17.260 14.750 ;
        RECT 14.310 13.220 14.600 14.630 ;
        RECT 14.940 13.760 15.110 14.090 ;
        RECT 15.325 14.060 16.365 14.230 ;
        RECT 15.325 13.620 16.365 13.790 ;
        RECT 16.580 13.760 16.750 14.090 ;
        RECT 17.090 13.220 17.260 14.630 ;
        RECT 14.310 13.100 17.260 13.220 ;
        RECT 14.430 13.050 17.260 13.100 ;
        RECT 17.820 14.720 20.560 14.790 ;
        RECT 21.140 14.720 23.880 14.790 ;
        RECT 17.820 14.620 20.690 14.720 ;
        RECT 17.820 13.210 17.990 14.620 ;
        RECT 18.330 13.750 18.500 14.080 ;
        RECT 18.670 14.050 19.710 14.220 ;
        RECT 18.670 13.610 19.710 13.780 ;
        RECT 19.880 13.750 20.050 14.080 ;
        RECT 20.390 13.210 20.690 14.620 ;
        RECT 17.820 13.070 20.690 13.210 ;
        RECT 21.010 14.620 23.880 14.720 ;
        RECT 21.010 13.210 21.310 14.620 ;
        RECT 21.650 13.750 21.820 14.080 ;
        RECT 21.990 14.050 23.030 14.220 ;
        RECT 21.990 13.610 23.030 13.780 ;
        RECT 23.200 13.750 23.370 14.080 ;
        RECT 23.710 13.210 23.880 14.620 ;
        RECT 21.010 13.070 23.880 13.210 ;
        RECT 17.820 13.040 20.560 13.070 ;
        RECT 21.140 13.040 23.880 13.070 ;
        RECT 24.440 14.750 27.270 14.800 ;
        RECT 24.440 14.630 27.390 14.750 ;
        RECT 24.440 13.220 24.610 14.630 ;
        RECT 24.950 13.760 25.120 14.090 ;
        RECT 25.335 14.060 26.375 14.230 ;
        RECT 25.335 13.620 26.375 13.790 ;
        RECT 26.590 13.760 26.760 14.090 ;
        RECT 27.100 13.220 27.390 14.630 ;
        RECT 24.440 13.100 27.390 13.220 ;
        RECT 24.440 13.050 27.270 13.100 ;
        RECT 14.430 12.650 17.260 12.700 ;
        RECT 14.310 12.530 17.260 12.650 ;
        RECT 14.310 11.120 14.600 12.530 ;
        RECT 14.940 11.660 15.110 11.990 ;
        RECT 15.325 11.960 16.365 12.130 ;
        RECT 15.325 11.520 16.365 11.690 ;
        RECT 16.580 11.660 16.750 11.990 ;
        RECT 17.090 11.120 17.260 12.530 ;
        RECT 14.310 11.000 17.260 11.120 ;
        RECT 14.430 10.950 17.260 11.000 ;
        RECT 17.820 12.620 20.560 12.690 ;
        RECT 21.140 12.620 23.880 12.690 ;
        RECT 17.820 12.520 20.690 12.620 ;
        RECT 17.820 11.110 17.990 12.520 ;
        RECT 18.330 11.650 18.500 11.980 ;
        RECT 18.670 11.950 19.710 12.120 ;
        RECT 18.670 11.510 19.710 11.680 ;
        RECT 19.880 11.650 20.050 11.980 ;
        RECT 20.390 11.110 20.690 12.520 ;
        RECT 17.820 10.970 20.690 11.110 ;
        RECT 21.010 12.520 23.880 12.620 ;
        RECT 21.010 11.110 21.310 12.520 ;
        RECT 21.650 11.650 21.820 11.980 ;
        RECT 21.990 11.950 23.030 12.120 ;
        RECT 21.990 11.510 23.030 11.680 ;
        RECT 23.200 11.650 23.370 11.980 ;
        RECT 23.710 11.110 23.880 12.520 ;
        RECT 21.010 10.970 23.880 11.110 ;
        RECT 17.820 10.940 20.560 10.970 ;
        RECT 21.140 10.940 23.880 10.970 ;
        RECT 24.440 12.650 27.270 12.700 ;
        RECT 24.440 12.530 27.390 12.650 ;
        RECT 24.440 11.120 24.610 12.530 ;
        RECT 24.950 11.660 25.120 11.990 ;
        RECT 25.335 11.960 26.375 12.130 ;
        RECT 25.335 11.520 26.375 11.690 ;
        RECT 26.590 11.660 26.760 11.990 ;
        RECT 27.100 11.120 27.390 12.530 ;
        RECT 24.440 11.000 27.390 11.120 ;
        RECT 24.440 10.950 27.270 11.000 ;
      LAYER mcon ;
        RECT 15.405 219.800 16.285 219.970 ;
        RECT 14.940 219.580 15.110 219.750 ;
        RECT 16.580 219.580 16.750 219.750 ;
        RECT 15.405 219.360 16.285 219.530 ;
        RECT 18.750 219.790 19.630 219.960 ;
        RECT 18.330 219.570 18.500 219.740 ;
        RECT 19.880 219.570 20.050 219.740 ;
        RECT 18.750 219.350 19.630 219.520 ;
        RECT 20.430 218.810 20.690 220.460 ;
        RECT 22.070 219.850 22.950 220.020 ;
        RECT 21.650 219.630 21.820 219.800 ;
        RECT 23.200 219.630 23.370 219.800 ;
        RECT 22.070 219.410 22.950 219.580 ;
        RECT 25.415 219.860 26.295 220.030 ;
        RECT 24.950 219.640 25.120 219.810 ;
        RECT 26.590 219.640 26.760 219.810 ;
        RECT 25.415 219.420 26.295 219.590 ;
        RECT 15.405 217.700 16.285 217.870 ;
        RECT 14.940 217.480 15.110 217.650 ;
        RECT 16.580 217.480 16.750 217.650 ;
        RECT 15.405 217.260 16.285 217.430 ;
        RECT 18.750 217.690 19.630 217.860 ;
        RECT 18.330 217.470 18.500 217.640 ;
        RECT 19.880 217.470 20.050 217.640 ;
        RECT 18.750 217.250 19.630 217.420 ;
        RECT 20.430 216.710 20.690 218.360 ;
        RECT 27.130 218.900 27.390 220.550 ;
        RECT 22.070 217.750 22.950 217.920 ;
        RECT 21.650 217.530 21.820 217.700 ;
        RECT 23.200 217.530 23.370 217.700 ;
        RECT 22.070 217.310 22.950 217.480 ;
        RECT 25.415 217.760 26.295 217.930 ;
        RECT 24.950 217.540 25.120 217.710 ;
        RECT 26.590 217.540 26.760 217.710 ;
        RECT 25.415 217.320 26.295 217.490 ;
        RECT 15.405 215.600 16.285 215.770 ;
        RECT 14.940 215.380 15.110 215.550 ;
        RECT 16.580 215.380 16.750 215.550 ;
        RECT 15.405 215.160 16.285 215.330 ;
        RECT 18.750 215.590 19.630 215.760 ;
        RECT 18.330 215.370 18.500 215.540 ;
        RECT 19.880 215.370 20.050 215.540 ;
        RECT 18.750 215.150 19.630 215.320 ;
        RECT 20.430 214.610 20.690 216.260 ;
        RECT 27.130 216.800 27.390 218.450 ;
        RECT 22.070 215.650 22.950 215.820 ;
        RECT 21.650 215.430 21.820 215.600 ;
        RECT 23.200 215.430 23.370 215.600 ;
        RECT 22.070 215.210 22.950 215.380 ;
        RECT 15.405 213.500 16.285 213.670 ;
        RECT 14.940 213.280 15.110 213.450 ;
        RECT 16.580 213.280 16.750 213.450 ;
        RECT 15.405 213.060 16.285 213.230 ;
        RECT 25.415 215.660 26.295 215.830 ;
        RECT 24.950 215.440 25.120 215.610 ;
        RECT 26.590 215.440 26.760 215.610 ;
        RECT 25.415 215.220 26.295 215.390 ;
        RECT 27.130 214.700 27.390 216.350 ;
        RECT 18.750 213.490 19.630 213.660 ;
        RECT 18.330 213.270 18.500 213.440 ;
        RECT 19.880 213.270 20.050 213.440 ;
        RECT 18.750 213.050 19.630 213.220 ;
        RECT 20.430 212.510 20.690 214.160 ;
        RECT 22.070 213.550 22.950 213.720 ;
        RECT 21.650 213.330 21.820 213.500 ;
        RECT 23.200 213.330 23.370 213.500 ;
        RECT 22.070 213.110 22.950 213.280 ;
        RECT 25.415 213.560 26.295 213.730 ;
        RECT 24.950 213.340 25.120 213.510 ;
        RECT 26.590 213.340 26.760 213.510 ;
        RECT 25.415 213.120 26.295 213.290 ;
        RECT 27.130 212.600 27.390 214.250 ;
        RECT 15.405 211.410 16.285 211.580 ;
        RECT 14.940 211.190 15.110 211.360 ;
        RECT 16.580 211.190 16.750 211.360 ;
        RECT 15.405 210.970 16.285 211.140 ;
        RECT 18.750 211.400 19.630 211.570 ;
        RECT 18.330 211.180 18.500 211.350 ;
        RECT 19.880 211.180 20.050 211.350 ;
        RECT 18.750 210.960 19.630 211.130 ;
        RECT 20.430 210.420 20.690 212.070 ;
        RECT 22.070 211.450 22.950 211.620 ;
        RECT 21.650 211.230 21.820 211.400 ;
        RECT 23.200 211.230 23.370 211.400 ;
        RECT 22.070 211.010 22.950 211.180 ;
        RECT 25.415 211.460 26.295 211.630 ;
        RECT 24.950 211.240 25.120 211.410 ;
        RECT 26.590 211.240 26.760 211.410 ;
        RECT 25.415 211.020 26.295 211.190 ;
        RECT 27.130 210.500 27.390 212.150 ;
        RECT 15.405 209.310 16.285 209.480 ;
        RECT 14.940 209.090 15.110 209.260 ;
        RECT 16.580 209.090 16.750 209.260 ;
        RECT 15.405 208.870 16.285 209.040 ;
        RECT 18.750 209.300 19.630 209.470 ;
        RECT 18.330 209.080 18.500 209.250 ;
        RECT 19.880 209.080 20.050 209.250 ;
        RECT 18.750 208.860 19.630 209.030 ;
        RECT 20.430 208.320 20.690 209.970 ;
        RECT 22.070 209.350 22.950 209.520 ;
        RECT 21.650 209.130 21.820 209.300 ;
        RECT 23.200 209.130 23.370 209.300 ;
        RECT 22.070 208.910 22.950 209.080 ;
        RECT 25.415 209.360 26.295 209.530 ;
        RECT 24.950 209.140 25.120 209.310 ;
        RECT 26.590 209.140 26.760 209.310 ;
        RECT 25.415 208.920 26.295 209.090 ;
        RECT 27.130 208.400 27.390 210.050 ;
        RECT 15.405 207.220 16.285 207.390 ;
        RECT 14.940 207.000 15.110 207.170 ;
        RECT 16.580 207.000 16.750 207.170 ;
        RECT 15.405 206.780 16.285 206.950 ;
        RECT 18.750 207.210 19.630 207.380 ;
        RECT 18.330 206.990 18.500 207.160 ;
        RECT 19.880 206.990 20.050 207.160 ;
        RECT 18.750 206.770 19.630 206.940 ;
        RECT 20.430 206.230 20.690 207.880 ;
        RECT 22.070 207.250 22.950 207.420 ;
        RECT 21.650 207.030 21.820 207.200 ;
        RECT 23.200 207.030 23.370 207.200 ;
        RECT 22.070 206.810 22.950 206.980 ;
        RECT 25.415 207.260 26.295 207.430 ;
        RECT 24.950 207.040 25.120 207.210 ;
        RECT 26.590 207.040 26.760 207.210 ;
        RECT 25.415 206.820 26.295 206.990 ;
        RECT 27.130 206.300 27.390 207.950 ;
        RECT 15.405 205.120 16.285 205.290 ;
        RECT 14.940 204.900 15.110 205.070 ;
        RECT 16.580 204.900 16.750 205.070 ;
        RECT 15.405 204.680 16.285 204.850 ;
        RECT 18.750 205.110 19.630 205.280 ;
        RECT 18.330 204.890 18.500 205.060 ;
        RECT 19.880 204.890 20.050 205.060 ;
        RECT 18.750 204.670 19.630 204.840 ;
        RECT 20.430 204.130 20.690 205.780 ;
        RECT 22.070 205.150 22.950 205.320 ;
        RECT 21.650 204.930 21.820 205.100 ;
        RECT 23.200 204.930 23.370 205.100 ;
        RECT 22.070 204.710 22.950 204.880 ;
        RECT 25.415 205.160 26.295 205.330 ;
        RECT 24.950 204.940 25.120 205.110 ;
        RECT 26.590 204.940 26.760 205.110 ;
        RECT 25.415 204.720 26.295 204.890 ;
        RECT 27.130 204.200 27.390 205.850 ;
        RECT 15.405 203.020 16.285 203.190 ;
        RECT 14.940 202.800 15.110 202.970 ;
        RECT 16.580 202.800 16.750 202.970 ;
        RECT 15.405 202.580 16.285 202.750 ;
        RECT 18.750 203.010 19.630 203.180 ;
        RECT 18.330 202.790 18.500 202.960 ;
        RECT 19.880 202.790 20.050 202.960 ;
        RECT 18.750 202.570 19.630 202.740 ;
        RECT 20.430 202.030 20.690 203.680 ;
        RECT 22.070 203.050 22.950 203.220 ;
        RECT 21.650 202.830 21.820 203.000 ;
        RECT 23.200 202.830 23.370 203.000 ;
        RECT 22.070 202.610 22.950 202.780 ;
        RECT 25.415 203.060 26.295 203.230 ;
        RECT 24.950 202.840 25.120 203.010 ;
        RECT 26.590 202.840 26.760 203.010 ;
        RECT 25.415 202.620 26.295 202.790 ;
        RECT 27.130 202.100 27.390 203.750 ;
        RECT 15.405 200.920 16.285 201.090 ;
        RECT 14.940 200.700 15.110 200.870 ;
        RECT 16.580 200.700 16.750 200.870 ;
        RECT 15.405 200.480 16.285 200.650 ;
        RECT 18.750 200.910 19.630 201.080 ;
        RECT 18.330 200.690 18.500 200.860 ;
        RECT 19.880 200.690 20.050 200.860 ;
        RECT 18.750 200.470 19.630 200.640 ;
        RECT 20.430 199.930 20.690 201.580 ;
        RECT 22.070 200.950 22.950 201.120 ;
        RECT 21.650 200.730 21.820 200.900 ;
        RECT 23.200 200.730 23.370 200.900 ;
        RECT 22.070 200.510 22.950 200.680 ;
        RECT 25.415 200.960 26.295 201.130 ;
        RECT 24.950 200.740 25.120 200.910 ;
        RECT 26.590 200.740 26.760 200.910 ;
        RECT 25.415 200.520 26.295 200.690 ;
        RECT 27.130 200.000 27.390 201.650 ;
        RECT 15.405 198.820 16.285 198.990 ;
        RECT 14.940 198.600 15.110 198.770 ;
        RECT 16.580 198.600 16.750 198.770 ;
        RECT 15.405 198.380 16.285 198.550 ;
        RECT 18.750 198.810 19.630 198.980 ;
        RECT 18.330 198.590 18.500 198.760 ;
        RECT 19.880 198.590 20.050 198.760 ;
        RECT 18.750 198.370 19.630 198.540 ;
        RECT 20.430 197.830 20.690 199.480 ;
        RECT 22.070 198.850 22.950 199.020 ;
        RECT 21.650 198.630 21.820 198.800 ;
        RECT 23.200 198.630 23.370 198.800 ;
        RECT 22.070 198.410 22.950 198.580 ;
        RECT 25.415 198.860 26.295 199.030 ;
        RECT 24.950 198.640 25.120 198.810 ;
        RECT 26.590 198.640 26.760 198.810 ;
        RECT 25.415 198.420 26.295 198.590 ;
        RECT 27.130 197.900 27.390 199.550 ;
        RECT 15.405 196.720 16.285 196.890 ;
        RECT 14.940 196.500 15.110 196.670 ;
        RECT 16.580 196.500 16.750 196.670 ;
        RECT 15.405 196.280 16.285 196.450 ;
        RECT 18.750 196.710 19.630 196.880 ;
        RECT 18.330 196.490 18.500 196.660 ;
        RECT 19.880 196.490 20.050 196.660 ;
        RECT 18.750 196.270 19.630 196.440 ;
        RECT 20.430 195.730 20.690 197.380 ;
        RECT 22.070 196.750 22.950 196.920 ;
        RECT 21.650 196.530 21.820 196.700 ;
        RECT 23.200 196.530 23.370 196.700 ;
        RECT 22.070 196.310 22.950 196.480 ;
        RECT 25.415 196.760 26.295 196.930 ;
        RECT 24.950 196.540 25.120 196.710 ;
        RECT 26.590 196.540 26.760 196.710 ;
        RECT 25.415 196.320 26.295 196.490 ;
        RECT 27.130 195.800 27.390 197.450 ;
        RECT 15.405 194.620 16.285 194.790 ;
        RECT 14.940 194.400 15.110 194.570 ;
        RECT 16.580 194.400 16.750 194.570 ;
        RECT 15.405 194.180 16.285 194.350 ;
        RECT 18.750 194.610 19.630 194.780 ;
        RECT 18.330 194.390 18.500 194.560 ;
        RECT 19.880 194.390 20.050 194.560 ;
        RECT 18.750 194.170 19.630 194.340 ;
        RECT 20.430 193.630 20.690 195.280 ;
        RECT 22.070 194.650 22.950 194.820 ;
        RECT 21.650 194.430 21.820 194.600 ;
        RECT 23.200 194.430 23.370 194.600 ;
        RECT 22.070 194.210 22.950 194.380 ;
        RECT 25.415 194.660 26.295 194.830 ;
        RECT 24.950 194.440 25.120 194.610 ;
        RECT 26.590 194.440 26.760 194.610 ;
        RECT 25.415 194.220 26.295 194.390 ;
        RECT 27.130 193.700 27.390 195.350 ;
        RECT 15.405 192.520 16.285 192.690 ;
        RECT 14.940 192.300 15.110 192.470 ;
        RECT 16.580 192.300 16.750 192.470 ;
        RECT 15.405 192.080 16.285 192.250 ;
        RECT 18.750 192.510 19.630 192.680 ;
        RECT 18.330 192.290 18.500 192.460 ;
        RECT 19.880 192.290 20.050 192.460 ;
        RECT 18.750 192.070 19.630 192.240 ;
        RECT 20.430 191.530 20.690 193.180 ;
        RECT 22.070 192.550 22.950 192.720 ;
        RECT 21.650 192.330 21.820 192.500 ;
        RECT 23.200 192.330 23.370 192.500 ;
        RECT 22.070 192.110 22.950 192.280 ;
        RECT 25.415 192.560 26.295 192.730 ;
        RECT 24.950 192.340 25.120 192.510 ;
        RECT 26.590 192.340 26.760 192.510 ;
        RECT 25.415 192.120 26.295 192.290 ;
        RECT 27.130 191.600 27.390 193.250 ;
        RECT 15.405 190.420 16.285 190.590 ;
        RECT 14.940 190.200 15.110 190.370 ;
        RECT 16.580 190.200 16.750 190.370 ;
        RECT 15.405 189.980 16.285 190.150 ;
        RECT 18.750 190.410 19.630 190.580 ;
        RECT 18.330 190.190 18.500 190.360 ;
        RECT 19.880 190.190 20.050 190.360 ;
        RECT 18.750 189.970 19.630 190.140 ;
        RECT 20.430 189.430 20.690 191.080 ;
        RECT 22.070 190.450 22.950 190.620 ;
        RECT 21.650 190.230 21.820 190.400 ;
        RECT 23.200 190.230 23.370 190.400 ;
        RECT 22.070 190.010 22.950 190.180 ;
        RECT 25.415 190.460 26.295 190.630 ;
        RECT 24.950 190.240 25.120 190.410 ;
        RECT 26.590 190.240 26.760 190.410 ;
        RECT 25.415 190.020 26.295 190.190 ;
        RECT 27.130 189.500 27.390 191.150 ;
        RECT 15.405 188.330 16.285 188.500 ;
        RECT 14.940 188.110 15.110 188.280 ;
        RECT 16.580 188.110 16.750 188.280 ;
        RECT 15.405 187.890 16.285 188.060 ;
        RECT 18.750 188.320 19.630 188.490 ;
        RECT 18.330 188.100 18.500 188.270 ;
        RECT 19.880 188.100 20.050 188.270 ;
        RECT 18.750 187.880 19.630 188.050 ;
        RECT 20.430 187.340 20.690 188.990 ;
        RECT 22.070 188.350 22.950 188.520 ;
        RECT 21.650 188.130 21.820 188.300 ;
        RECT 23.200 188.130 23.370 188.300 ;
        RECT 22.070 187.910 22.950 188.080 ;
        RECT 25.415 188.360 26.295 188.530 ;
        RECT 24.950 188.140 25.120 188.310 ;
        RECT 26.590 188.140 26.760 188.310 ;
        RECT 25.415 187.920 26.295 188.090 ;
        RECT 27.130 187.400 27.390 189.050 ;
        RECT 15.405 186.240 16.285 186.410 ;
        RECT 14.940 186.020 15.110 186.190 ;
        RECT 16.580 186.020 16.750 186.190 ;
        RECT 15.405 185.800 16.285 185.970 ;
        RECT 18.750 186.230 19.630 186.400 ;
        RECT 18.330 186.010 18.500 186.180 ;
        RECT 19.880 186.010 20.050 186.180 ;
        RECT 18.750 185.790 19.630 185.960 ;
        RECT 20.430 185.250 20.690 186.900 ;
        RECT 22.070 186.250 22.950 186.420 ;
        RECT 21.650 186.030 21.820 186.200 ;
        RECT 23.200 186.030 23.370 186.200 ;
        RECT 22.070 185.810 22.950 185.980 ;
        RECT 25.415 186.260 26.295 186.430 ;
        RECT 24.950 186.040 25.120 186.210 ;
        RECT 26.590 186.040 26.760 186.210 ;
        RECT 25.415 185.820 26.295 185.990 ;
        RECT 27.130 185.300 27.390 186.950 ;
        RECT 15.405 184.140 16.285 184.310 ;
        RECT 14.940 183.920 15.110 184.090 ;
        RECT 16.580 183.920 16.750 184.090 ;
        RECT 15.405 183.700 16.285 183.870 ;
        RECT 18.750 184.130 19.630 184.300 ;
        RECT 18.330 183.910 18.500 184.080 ;
        RECT 19.880 183.910 20.050 184.080 ;
        RECT 18.750 183.690 19.630 183.860 ;
        RECT 20.430 183.150 20.690 184.800 ;
        RECT 22.070 184.150 22.950 184.320 ;
        RECT 21.650 183.930 21.820 184.100 ;
        RECT 23.200 183.930 23.370 184.100 ;
        RECT 22.070 183.710 22.950 183.880 ;
        RECT 25.415 184.160 26.295 184.330 ;
        RECT 24.950 183.940 25.120 184.110 ;
        RECT 26.590 183.940 26.760 184.110 ;
        RECT 25.415 183.720 26.295 183.890 ;
        RECT 27.130 183.200 27.390 184.850 ;
        RECT 15.405 182.050 16.285 182.220 ;
        RECT 14.940 181.830 15.110 182.000 ;
        RECT 16.580 181.830 16.750 182.000 ;
        RECT 15.405 181.610 16.285 181.780 ;
        RECT 18.750 182.040 19.630 182.210 ;
        RECT 18.330 181.820 18.500 181.990 ;
        RECT 19.880 181.820 20.050 181.990 ;
        RECT 18.750 181.600 19.630 181.770 ;
        RECT 20.430 181.060 20.690 182.710 ;
        RECT 22.070 182.050 22.950 182.220 ;
        RECT 21.650 181.830 21.820 182.000 ;
        RECT 23.200 181.830 23.370 182.000 ;
        RECT 22.070 181.610 22.950 181.780 ;
        RECT 25.415 182.060 26.295 182.230 ;
        RECT 24.950 181.840 25.120 182.010 ;
        RECT 26.590 181.840 26.760 182.010 ;
        RECT 25.415 181.620 26.295 181.790 ;
        RECT 27.130 181.100 27.390 182.750 ;
        RECT 15.405 179.960 16.285 180.130 ;
        RECT 14.940 179.740 15.110 179.910 ;
        RECT 16.580 179.740 16.750 179.910 ;
        RECT 15.405 179.520 16.285 179.690 ;
        RECT 18.750 179.950 19.630 180.120 ;
        RECT 18.330 179.730 18.500 179.900 ;
        RECT 19.880 179.730 20.050 179.900 ;
        RECT 18.750 179.510 19.630 179.680 ;
        RECT 20.430 178.970 20.690 180.620 ;
        RECT 22.070 179.950 22.950 180.120 ;
        RECT 21.650 179.730 21.820 179.900 ;
        RECT 23.200 179.730 23.370 179.900 ;
        RECT 22.070 179.510 22.950 179.680 ;
        RECT 25.415 179.960 26.295 180.130 ;
        RECT 24.950 179.740 25.120 179.910 ;
        RECT 26.590 179.740 26.760 179.910 ;
        RECT 25.415 179.520 26.295 179.690 ;
        RECT 27.130 179.000 27.390 180.650 ;
        RECT 15.405 177.860 16.285 178.030 ;
        RECT 14.940 177.640 15.110 177.810 ;
        RECT 16.580 177.640 16.750 177.810 ;
        RECT 15.405 177.420 16.285 177.590 ;
        RECT 18.750 177.850 19.630 178.020 ;
        RECT 18.330 177.630 18.500 177.800 ;
        RECT 19.880 177.630 20.050 177.800 ;
        RECT 18.750 177.410 19.630 177.580 ;
        RECT 20.430 176.870 20.690 178.520 ;
        RECT 22.070 177.850 22.950 178.020 ;
        RECT 21.650 177.630 21.820 177.800 ;
        RECT 23.200 177.630 23.370 177.800 ;
        RECT 22.070 177.410 22.950 177.580 ;
        RECT 25.415 177.860 26.295 178.030 ;
        RECT 24.950 177.640 25.120 177.810 ;
        RECT 26.590 177.640 26.760 177.810 ;
        RECT 25.415 177.420 26.295 177.590 ;
        RECT 27.130 176.900 27.390 178.550 ;
        RECT 15.405 175.760 16.285 175.930 ;
        RECT 14.940 175.540 15.110 175.710 ;
        RECT 16.580 175.540 16.750 175.710 ;
        RECT 15.405 175.320 16.285 175.490 ;
        RECT 18.750 175.750 19.630 175.920 ;
        RECT 18.330 175.530 18.500 175.700 ;
        RECT 19.880 175.530 20.050 175.700 ;
        RECT 18.750 175.310 19.630 175.480 ;
        RECT 20.430 174.770 20.690 176.420 ;
        RECT 22.070 175.750 22.950 175.920 ;
        RECT 21.650 175.530 21.820 175.700 ;
        RECT 23.200 175.530 23.370 175.700 ;
        RECT 22.070 175.310 22.950 175.480 ;
        RECT 25.415 175.760 26.295 175.930 ;
        RECT 24.950 175.540 25.120 175.710 ;
        RECT 26.590 175.540 26.760 175.710 ;
        RECT 25.415 175.320 26.295 175.490 ;
        RECT 27.130 174.800 27.390 176.450 ;
        RECT 15.405 173.660 16.285 173.830 ;
        RECT 14.940 173.440 15.110 173.610 ;
        RECT 16.580 173.440 16.750 173.610 ;
        RECT 15.405 173.220 16.285 173.390 ;
        RECT 18.750 173.650 19.630 173.820 ;
        RECT 18.330 173.430 18.500 173.600 ;
        RECT 19.880 173.430 20.050 173.600 ;
        RECT 18.750 173.210 19.630 173.380 ;
        RECT 20.430 172.670 20.690 174.320 ;
        RECT 22.070 173.650 22.950 173.820 ;
        RECT 21.650 173.430 21.820 173.600 ;
        RECT 23.200 173.430 23.370 173.600 ;
        RECT 22.070 173.210 22.950 173.380 ;
        RECT 25.415 173.660 26.295 173.830 ;
        RECT 24.950 173.440 25.120 173.610 ;
        RECT 26.590 173.440 26.760 173.610 ;
        RECT 25.415 173.220 26.295 173.390 ;
        RECT 27.130 172.700 27.390 174.350 ;
        RECT 15.405 171.560 16.285 171.730 ;
        RECT 14.940 171.340 15.110 171.510 ;
        RECT 16.580 171.340 16.750 171.510 ;
        RECT 15.405 171.120 16.285 171.290 ;
        RECT 18.750 171.550 19.630 171.720 ;
        RECT 18.330 171.330 18.500 171.500 ;
        RECT 19.880 171.330 20.050 171.500 ;
        RECT 18.750 171.110 19.630 171.280 ;
        RECT 20.430 170.570 20.690 172.220 ;
        RECT 22.070 171.550 22.950 171.720 ;
        RECT 21.650 171.330 21.820 171.500 ;
        RECT 23.200 171.330 23.370 171.500 ;
        RECT 22.070 171.110 22.950 171.280 ;
        RECT 25.415 171.560 26.295 171.730 ;
        RECT 24.950 171.340 25.120 171.510 ;
        RECT 26.590 171.340 26.760 171.510 ;
        RECT 25.415 171.120 26.295 171.290 ;
        RECT 27.130 170.600 27.390 172.250 ;
        RECT 15.405 169.460 16.285 169.630 ;
        RECT 14.940 169.240 15.110 169.410 ;
        RECT 16.580 169.240 16.750 169.410 ;
        RECT 15.405 169.020 16.285 169.190 ;
        RECT 18.750 169.450 19.630 169.620 ;
        RECT 18.330 169.230 18.500 169.400 ;
        RECT 19.880 169.230 20.050 169.400 ;
        RECT 18.750 169.010 19.630 169.180 ;
        RECT 20.430 168.470 20.690 170.120 ;
        RECT 22.070 169.450 22.950 169.620 ;
        RECT 21.650 169.230 21.820 169.400 ;
        RECT 23.200 169.230 23.370 169.400 ;
        RECT 22.070 169.010 22.950 169.180 ;
        RECT 25.415 169.460 26.295 169.630 ;
        RECT 24.950 169.240 25.120 169.410 ;
        RECT 26.590 169.240 26.760 169.410 ;
        RECT 25.415 169.020 26.295 169.190 ;
        RECT 27.130 168.500 27.390 170.150 ;
        RECT 15.405 167.360 16.285 167.530 ;
        RECT 14.940 167.140 15.110 167.310 ;
        RECT 16.580 167.140 16.750 167.310 ;
        RECT 15.405 166.920 16.285 167.090 ;
        RECT 18.750 167.350 19.630 167.520 ;
        RECT 18.330 167.130 18.500 167.300 ;
        RECT 19.880 167.130 20.050 167.300 ;
        RECT 18.750 166.910 19.630 167.080 ;
        RECT 20.430 166.370 20.690 168.020 ;
        RECT 22.070 167.350 22.950 167.520 ;
        RECT 21.650 167.130 21.820 167.300 ;
        RECT 23.200 167.130 23.370 167.300 ;
        RECT 22.070 166.910 22.950 167.080 ;
        RECT 25.415 167.360 26.295 167.530 ;
        RECT 24.950 167.140 25.120 167.310 ;
        RECT 26.590 167.140 26.760 167.310 ;
        RECT 25.415 166.920 26.295 167.090 ;
        RECT 27.130 166.400 27.390 168.050 ;
        RECT 15.405 165.260 16.285 165.430 ;
        RECT 14.940 165.040 15.110 165.210 ;
        RECT 16.580 165.040 16.750 165.210 ;
        RECT 15.405 164.820 16.285 164.990 ;
        RECT 18.750 165.250 19.630 165.420 ;
        RECT 18.330 165.030 18.500 165.200 ;
        RECT 19.880 165.030 20.050 165.200 ;
        RECT 18.750 164.810 19.630 164.980 ;
        RECT 20.430 164.270 20.690 165.920 ;
        RECT 22.070 165.250 22.950 165.420 ;
        RECT 21.650 165.030 21.820 165.200 ;
        RECT 23.200 165.030 23.370 165.200 ;
        RECT 22.070 164.810 22.950 164.980 ;
        RECT 25.415 165.260 26.295 165.430 ;
        RECT 24.950 165.040 25.120 165.210 ;
        RECT 26.590 165.040 26.760 165.210 ;
        RECT 25.415 164.820 26.295 164.990 ;
        RECT 27.130 164.300 27.390 165.950 ;
        RECT 15.405 163.160 16.285 163.330 ;
        RECT 14.940 162.940 15.110 163.110 ;
        RECT 16.580 162.940 16.750 163.110 ;
        RECT 15.405 162.720 16.285 162.890 ;
        RECT 18.750 163.150 19.630 163.320 ;
        RECT 18.330 162.930 18.500 163.100 ;
        RECT 19.880 162.930 20.050 163.100 ;
        RECT 18.750 162.710 19.630 162.880 ;
        RECT 20.430 162.170 20.690 163.820 ;
        RECT 22.070 163.150 22.950 163.320 ;
        RECT 21.650 162.930 21.820 163.100 ;
        RECT 23.200 162.930 23.370 163.100 ;
        RECT 22.070 162.710 22.950 162.880 ;
        RECT 25.415 163.160 26.295 163.330 ;
        RECT 24.950 162.940 25.120 163.110 ;
        RECT 26.590 162.940 26.760 163.110 ;
        RECT 25.415 162.720 26.295 162.890 ;
        RECT 27.130 162.200 27.390 163.850 ;
        RECT 15.405 161.060 16.285 161.230 ;
        RECT 14.940 160.840 15.110 161.010 ;
        RECT 16.580 160.840 16.750 161.010 ;
        RECT 15.405 160.620 16.285 160.790 ;
        RECT 18.750 161.050 19.630 161.220 ;
        RECT 18.330 160.830 18.500 161.000 ;
        RECT 19.880 160.830 20.050 161.000 ;
        RECT 18.750 160.610 19.630 160.780 ;
        RECT 20.430 160.070 20.690 161.720 ;
        RECT 22.070 161.050 22.950 161.220 ;
        RECT 21.650 160.830 21.820 161.000 ;
        RECT 23.200 160.830 23.370 161.000 ;
        RECT 22.070 160.610 22.950 160.780 ;
        RECT 25.415 161.060 26.295 161.230 ;
        RECT 24.950 160.840 25.120 161.010 ;
        RECT 26.590 160.840 26.760 161.010 ;
        RECT 25.415 160.620 26.295 160.790 ;
        RECT 27.130 160.100 27.390 161.750 ;
        RECT 15.405 158.960 16.285 159.130 ;
        RECT 14.940 158.740 15.110 158.910 ;
        RECT 16.580 158.740 16.750 158.910 ;
        RECT 15.405 158.520 16.285 158.690 ;
        RECT 18.750 158.950 19.630 159.120 ;
        RECT 18.330 158.730 18.500 158.900 ;
        RECT 19.880 158.730 20.050 158.900 ;
        RECT 18.750 158.510 19.630 158.680 ;
        RECT 20.430 157.970 20.690 159.620 ;
        RECT 22.070 158.950 22.950 159.120 ;
        RECT 21.650 158.730 21.820 158.900 ;
        RECT 23.200 158.730 23.370 158.900 ;
        RECT 22.070 158.510 22.950 158.680 ;
        RECT 25.415 158.960 26.295 159.130 ;
        RECT 24.950 158.740 25.120 158.910 ;
        RECT 26.590 158.740 26.760 158.910 ;
        RECT 25.415 158.520 26.295 158.690 ;
        RECT 27.130 158.000 27.390 159.650 ;
        RECT 15.405 156.860 16.285 157.030 ;
        RECT 14.940 156.640 15.110 156.810 ;
        RECT 16.580 156.640 16.750 156.810 ;
        RECT 15.405 156.420 16.285 156.590 ;
        RECT 18.750 156.850 19.630 157.020 ;
        RECT 18.330 156.630 18.500 156.800 ;
        RECT 19.880 156.630 20.050 156.800 ;
        RECT 18.750 156.410 19.630 156.580 ;
        RECT 20.430 155.870 20.690 157.520 ;
        RECT 22.070 156.850 22.950 157.020 ;
        RECT 21.650 156.630 21.820 156.800 ;
        RECT 23.200 156.630 23.370 156.800 ;
        RECT 22.070 156.410 22.950 156.580 ;
        RECT 25.415 156.860 26.295 157.030 ;
        RECT 24.950 156.640 25.120 156.810 ;
        RECT 26.590 156.640 26.760 156.810 ;
        RECT 25.415 156.420 26.295 156.590 ;
        RECT 27.130 155.900 27.390 157.550 ;
        RECT 15.405 154.760 16.285 154.930 ;
        RECT 14.940 154.540 15.110 154.710 ;
        RECT 16.580 154.540 16.750 154.710 ;
        RECT 15.405 154.320 16.285 154.490 ;
        RECT 18.750 154.750 19.630 154.920 ;
        RECT 18.330 154.530 18.500 154.700 ;
        RECT 19.880 154.530 20.050 154.700 ;
        RECT 18.750 154.310 19.630 154.480 ;
        RECT 20.430 153.770 20.690 155.420 ;
        RECT 22.070 154.750 22.950 154.920 ;
        RECT 21.650 154.530 21.820 154.700 ;
        RECT 23.200 154.530 23.370 154.700 ;
        RECT 22.070 154.310 22.950 154.480 ;
        RECT 25.415 154.760 26.295 154.930 ;
        RECT 24.950 154.540 25.120 154.710 ;
        RECT 26.590 154.540 26.760 154.710 ;
        RECT 25.415 154.320 26.295 154.490 ;
        RECT 27.130 153.800 27.390 155.450 ;
        RECT 15.405 152.660 16.285 152.830 ;
        RECT 14.940 152.440 15.110 152.610 ;
        RECT 16.580 152.440 16.750 152.610 ;
        RECT 15.405 152.220 16.285 152.390 ;
        RECT 18.750 152.650 19.630 152.820 ;
        RECT 18.330 152.430 18.500 152.600 ;
        RECT 19.880 152.430 20.050 152.600 ;
        RECT 18.750 152.210 19.630 152.380 ;
        RECT 20.430 151.670 20.690 153.320 ;
        RECT 22.070 152.650 22.950 152.820 ;
        RECT 21.650 152.430 21.820 152.600 ;
        RECT 23.200 152.430 23.370 152.600 ;
        RECT 22.070 152.210 22.950 152.380 ;
        RECT 25.415 152.660 26.295 152.830 ;
        RECT 24.950 152.440 25.120 152.610 ;
        RECT 26.590 152.440 26.760 152.610 ;
        RECT 25.415 152.220 26.295 152.390 ;
        RECT 27.130 151.700 27.390 153.350 ;
        RECT 15.405 150.560 16.285 150.730 ;
        RECT 14.940 150.340 15.110 150.510 ;
        RECT 16.580 150.340 16.750 150.510 ;
        RECT 15.405 150.120 16.285 150.290 ;
        RECT 18.750 150.550 19.630 150.720 ;
        RECT 18.330 150.330 18.500 150.500 ;
        RECT 19.880 150.330 20.050 150.500 ;
        RECT 18.750 150.110 19.630 150.280 ;
        RECT 20.430 149.570 20.690 151.220 ;
        RECT 22.070 150.550 22.950 150.720 ;
        RECT 21.650 150.330 21.820 150.500 ;
        RECT 23.200 150.330 23.370 150.500 ;
        RECT 22.070 150.110 22.950 150.280 ;
        RECT 25.415 150.560 26.295 150.730 ;
        RECT 24.950 150.340 25.120 150.510 ;
        RECT 26.590 150.340 26.760 150.510 ;
        RECT 25.415 150.120 26.295 150.290 ;
        RECT 27.130 149.600 27.390 151.250 ;
        RECT 15.405 148.460 16.285 148.630 ;
        RECT 14.940 148.240 15.110 148.410 ;
        RECT 16.580 148.240 16.750 148.410 ;
        RECT 15.405 148.020 16.285 148.190 ;
        RECT 18.750 148.450 19.630 148.620 ;
        RECT 18.330 148.230 18.500 148.400 ;
        RECT 19.880 148.230 20.050 148.400 ;
        RECT 18.750 148.010 19.630 148.180 ;
        RECT 20.430 147.470 20.690 149.120 ;
        RECT 22.070 148.450 22.950 148.620 ;
        RECT 21.650 148.230 21.820 148.400 ;
        RECT 23.200 148.230 23.370 148.400 ;
        RECT 22.070 148.010 22.950 148.180 ;
        RECT 25.415 148.460 26.295 148.630 ;
        RECT 24.950 148.240 25.120 148.410 ;
        RECT 26.590 148.240 26.760 148.410 ;
        RECT 25.415 148.020 26.295 148.190 ;
        RECT 27.130 147.500 27.390 149.150 ;
        RECT 15.405 146.360 16.285 146.530 ;
        RECT 14.940 146.140 15.110 146.310 ;
        RECT 16.580 146.140 16.750 146.310 ;
        RECT 15.405 145.920 16.285 146.090 ;
        RECT 18.750 146.350 19.630 146.520 ;
        RECT 18.330 146.130 18.500 146.300 ;
        RECT 19.880 146.130 20.050 146.300 ;
        RECT 18.750 145.910 19.630 146.080 ;
        RECT 20.430 145.370 20.690 147.020 ;
        RECT 22.070 146.350 22.950 146.520 ;
        RECT 21.650 146.130 21.820 146.300 ;
        RECT 23.200 146.130 23.370 146.300 ;
        RECT 22.070 145.910 22.950 146.080 ;
        RECT 25.415 146.360 26.295 146.530 ;
        RECT 24.950 146.140 25.120 146.310 ;
        RECT 26.590 146.140 26.760 146.310 ;
        RECT 25.415 145.920 26.295 146.090 ;
        RECT 27.130 145.400 27.390 147.050 ;
        RECT 15.405 144.260 16.285 144.430 ;
        RECT 14.940 144.040 15.110 144.210 ;
        RECT 16.580 144.040 16.750 144.210 ;
        RECT 15.405 143.820 16.285 143.990 ;
        RECT 18.750 144.250 19.630 144.420 ;
        RECT 18.330 144.030 18.500 144.200 ;
        RECT 19.880 144.030 20.050 144.200 ;
        RECT 18.750 143.810 19.630 143.980 ;
        RECT 20.430 143.270 20.690 144.920 ;
        RECT 22.070 144.250 22.950 144.420 ;
        RECT 21.650 144.030 21.820 144.200 ;
        RECT 23.200 144.030 23.370 144.200 ;
        RECT 22.070 143.810 22.950 143.980 ;
        RECT 25.415 144.260 26.295 144.430 ;
        RECT 24.950 144.040 25.120 144.210 ;
        RECT 26.590 144.040 26.760 144.210 ;
        RECT 25.415 143.820 26.295 143.990 ;
        RECT 27.130 143.300 27.390 144.950 ;
        RECT 15.405 142.160 16.285 142.330 ;
        RECT 14.940 141.940 15.110 142.110 ;
        RECT 16.580 141.940 16.750 142.110 ;
        RECT 15.405 141.720 16.285 141.890 ;
        RECT 18.750 142.150 19.630 142.320 ;
        RECT 18.330 141.930 18.500 142.100 ;
        RECT 19.880 141.930 20.050 142.100 ;
        RECT 18.750 141.710 19.630 141.880 ;
        RECT 20.430 141.170 20.690 142.820 ;
        RECT 22.070 142.150 22.950 142.320 ;
        RECT 21.650 141.930 21.820 142.100 ;
        RECT 23.200 141.930 23.370 142.100 ;
        RECT 22.070 141.710 22.950 141.880 ;
        RECT 25.415 142.160 26.295 142.330 ;
        RECT 24.950 141.940 25.120 142.110 ;
        RECT 26.590 141.940 26.760 142.110 ;
        RECT 25.415 141.720 26.295 141.890 ;
        RECT 27.130 141.200 27.390 142.850 ;
        RECT 15.405 140.060 16.285 140.230 ;
        RECT 14.940 139.840 15.110 140.010 ;
        RECT 16.580 139.840 16.750 140.010 ;
        RECT 15.405 139.620 16.285 139.790 ;
        RECT 18.750 140.050 19.630 140.220 ;
        RECT 18.330 139.830 18.500 140.000 ;
        RECT 19.880 139.830 20.050 140.000 ;
        RECT 18.750 139.610 19.630 139.780 ;
        RECT 20.430 139.070 20.690 140.720 ;
        RECT 22.070 140.050 22.950 140.220 ;
        RECT 21.650 139.830 21.820 140.000 ;
        RECT 23.200 139.830 23.370 140.000 ;
        RECT 22.070 139.610 22.950 139.780 ;
        RECT 25.415 140.060 26.295 140.230 ;
        RECT 24.950 139.840 25.120 140.010 ;
        RECT 26.590 139.840 26.760 140.010 ;
        RECT 25.415 139.620 26.295 139.790 ;
        RECT 27.130 139.100 27.390 140.750 ;
        RECT 15.405 137.960 16.285 138.130 ;
        RECT 14.940 137.740 15.110 137.910 ;
        RECT 16.580 137.740 16.750 137.910 ;
        RECT 15.405 137.520 16.285 137.690 ;
        RECT 18.750 137.950 19.630 138.120 ;
        RECT 18.330 137.730 18.500 137.900 ;
        RECT 19.880 137.730 20.050 137.900 ;
        RECT 18.750 137.510 19.630 137.680 ;
        RECT 20.430 136.970 20.690 138.620 ;
        RECT 22.070 137.950 22.950 138.120 ;
        RECT 21.650 137.730 21.820 137.900 ;
        RECT 23.200 137.730 23.370 137.900 ;
        RECT 22.070 137.510 22.950 137.680 ;
        RECT 25.415 137.960 26.295 138.130 ;
        RECT 24.950 137.740 25.120 137.910 ;
        RECT 26.590 137.740 26.760 137.910 ;
        RECT 25.415 137.520 26.295 137.690 ;
        RECT 27.130 137.000 27.390 138.650 ;
        RECT 15.405 135.860 16.285 136.030 ;
        RECT 14.940 135.640 15.110 135.810 ;
        RECT 16.580 135.640 16.750 135.810 ;
        RECT 15.405 135.420 16.285 135.590 ;
        RECT 18.750 135.850 19.630 136.020 ;
        RECT 18.330 135.630 18.500 135.800 ;
        RECT 19.880 135.630 20.050 135.800 ;
        RECT 18.750 135.410 19.630 135.580 ;
        RECT 20.430 134.870 20.690 136.520 ;
        RECT 22.070 135.850 22.950 136.020 ;
        RECT 21.650 135.630 21.820 135.800 ;
        RECT 23.200 135.630 23.370 135.800 ;
        RECT 22.070 135.410 22.950 135.580 ;
        RECT 25.415 135.860 26.295 136.030 ;
        RECT 24.950 135.640 25.120 135.810 ;
        RECT 26.590 135.640 26.760 135.810 ;
        RECT 25.415 135.420 26.295 135.590 ;
        RECT 27.130 134.900 27.390 136.550 ;
        RECT 15.405 133.760 16.285 133.930 ;
        RECT 14.940 133.540 15.110 133.710 ;
        RECT 16.580 133.540 16.750 133.710 ;
        RECT 15.405 133.320 16.285 133.490 ;
        RECT 18.750 133.750 19.630 133.920 ;
        RECT 18.330 133.530 18.500 133.700 ;
        RECT 19.880 133.530 20.050 133.700 ;
        RECT 18.750 133.310 19.630 133.480 ;
        RECT 20.430 132.770 20.690 134.420 ;
        RECT 22.070 133.750 22.950 133.920 ;
        RECT 21.650 133.530 21.820 133.700 ;
        RECT 23.200 133.530 23.370 133.700 ;
        RECT 22.070 133.310 22.950 133.480 ;
        RECT 25.415 133.760 26.295 133.930 ;
        RECT 24.950 133.540 25.120 133.710 ;
        RECT 26.590 133.540 26.760 133.710 ;
        RECT 25.415 133.320 26.295 133.490 ;
        RECT 27.130 132.800 27.390 134.450 ;
        RECT 15.405 131.660 16.285 131.830 ;
        RECT 14.940 131.440 15.110 131.610 ;
        RECT 16.580 131.440 16.750 131.610 ;
        RECT 15.405 131.220 16.285 131.390 ;
        RECT 18.750 131.650 19.630 131.820 ;
        RECT 18.330 131.430 18.500 131.600 ;
        RECT 19.880 131.430 20.050 131.600 ;
        RECT 18.750 131.210 19.630 131.380 ;
        RECT 20.430 130.670 20.690 132.320 ;
        RECT 22.070 131.650 22.950 131.820 ;
        RECT 21.650 131.430 21.820 131.600 ;
        RECT 23.200 131.430 23.370 131.600 ;
        RECT 22.070 131.210 22.950 131.380 ;
        RECT 25.415 131.660 26.295 131.830 ;
        RECT 24.950 131.440 25.120 131.610 ;
        RECT 26.590 131.440 26.760 131.610 ;
        RECT 25.415 131.220 26.295 131.390 ;
        RECT 27.130 130.700 27.390 132.350 ;
        RECT 15.405 129.560 16.285 129.730 ;
        RECT 14.940 129.340 15.110 129.510 ;
        RECT 16.580 129.340 16.750 129.510 ;
        RECT 15.405 129.120 16.285 129.290 ;
        RECT 18.750 129.550 19.630 129.720 ;
        RECT 18.330 129.330 18.500 129.500 ;
        RECT 19.880 129.330 20.050 129.500 ;
        RECT 18.750 129.110 19.630 129.280 ;
        RECT 20.430 128.570 20.690 130.220 ;
        RECT 22.070 129.550 22.950 129.720 ;
        RECT 21.650 129.330 21.820 129.500 ;
        RECT 23.200 129.330 23.370 129.500 ;
        RECT 22.070 129.110 22.950 129.280 ;
        RECT 25.415 129.560 26.295 129.730 ;
        RECT 24.950 129.340 25.120 129.510 ;
        RECT 26.590 129.340 26.760 129.510 ;
        RECT 25.415 129.120 26.295 129.290 ;
        RECT 27.130 128.600 27.390 130.250 ;
        RECT 15.405 127.460 16.285 127.630 ;
        RECT 14.940 127.240 15.110 127.410 ;
        RECT 16.580 127.240 16.750 127.410 ;
        RECT 15.405 127.020 16.285 127.190 ;
        RECT 18.750 127.450 19.630 127.620 ;
        RECT 18.330 127.230 18.500 127.400 ;
        RECT 19.880 127.230 20.050 127.400 ;
        RECT 18.750 127.010 19.630 127.180 ;
        RECT 20.430 126.470 20.690 128.120 ;
        RECT 22.070 127.450 22.950 127.620 ;
        RECT 21.650 127.230 21.820 127.400 ;
        RECT 23.200 127.230 23.370 127.400 ;
        RECT 22.070 127.010 22.950 127.180 ;
        RECT 25.415 127.460 26.295 127.630 ;
        RECT 24.950 127.240 25.120 127.410 ;
        RECT 26.590 127.240 26.760 127.410 ;
        RECT 25.415 127.020 26.295 127.190 ;
        RECT 27.130 126.500 27.390 128.150 ;
        RECT 15.405 125.360 16.285 125.530 ;
        RECT 14.940 125.140 15.110 125.310 ;
        RECT 16.580 125.140 16.750 125.310 ;
        RECT 15.405 124.920 16.285 125.090 ;
        RECT 18.750 125.350 19.630 125.520 ;
        RECT 18.330 125.130 18.500 125.300 ;
        RECT 19.880 125.130 20.050 125.300 ;
        RECT 18.750 124.910 19.630 125.080 ;
        RECT 20.430 124.370 20.690 126.020 ;
        RECT 22.070 125.350 22.950 125.520 ;
        RECT 21.650 125.130 21.820 125.300 ;
        RECT 23.200 125.130 23.370 125.300 ;
        RECT 22.070 124.910 22.950 125.080 ;
        RECT 25.415 125.360 26.295 125.530 ;
        RECT 24.950 125.140 25.120 125.310 ;
        RECT 26.590 125.140 26.760 125.310 ;
        RECT 25.415 124.920 26.295 125.090 ;
        RECT 27.130 124.400 27.390 126.050 ;
        RECT 15.405 123.260 16.285 123.430 ;
        RECT 14.940 123.040 15.110 123.210 ;
        RECT 16.580 123.040 16.750 123.210 ;
        RECT 15.405 122.820 16.285 122.990 ;
        RECT 18.750 123.250 19.630 123.420 ;
        RECT 18.330 123.030 18.500 123.200 ;
        RECT 19.880 123.030 20.050 123.200 ;
        RECT 18.750 122.810 19.630 122.980 ;
        RECT 20.430 122.270 20.690 123.920 ;
        RECT 22.070 123.250 22.950 123.420 ;
        RECT 21.650 123.030 21.820 123.200 ;
        RECT 23.200 123.030 23.370 123.200 ;
        RECT 22.070 122.810 22.950 122.980 ;
        RECT 25.415 123.260 26.295 123.430 ;
        RECT 24.950 123.040 25.120 123.210 ;
        RECT 26.590 123.040 26.760 123.210 ;
        RECT 25.415 122.820 26.295 122.990 ;
        RECT 27.130 122.300 27.390 123.950 ;
        RECT 15.405 121.160 16.285 121.330 ;
        RECT 14.940 120.940 15.110 121.110 ;
        RECT 16.580 120.940 16.750 121.110 ;
        RECT 15.405 120.720 16.285 120.890 ;
        RECT 18.750 121.150 19.630 121.320 ;
        RECT 18.330 120.930 18.500 121.100 ;
        RECT 19.880 120.930 20.050 121.100 ;
        RECT 18.750 120.710 19.630 120.880 ;
        RECT 20.430 120.170 20.690 121.820 ;
        RECT 22.070 121.150 22.950 121.320 ;
        RECT 21.650 120.930 21.820 121.100 ;
        RECT 23.200 120.930 23.370 121.100 ;
        RECT 22.070 120.710 22.950 120.880 ;
        RECT 25.415 121.160 26.295 121.330 ;
        RECT 24.950 120.940 25.120 121.110 ;
        RECT 26.590 120.940 26.760 121.110 ;
        RECT 25.415 120.720 26.295 120.890 ;
        RECT 27.130 120.200 27.390 121.850 ;
        RECT 15.405 119.060 16.285 119.230 ;
        RECT 14.940 118.840 15.110 119.010 ;
        RECT 16.580 118.840 16.750 119.010 ;
        RECT 15.405 118.620 16.285 118.790 ;
        RECT 18.750 119.050 19.630 119.220 ;
        RECT 18.330 118.830 18.500 119.000 ;
        RECT 19.880 118.830 20.050 119.000 ;
        RECT 18.750 118.610 19.630 118.780 ;
        RECT 20.430 118.070 20.690 119.720 ;
        RECT 22.070 119.050 22.950 119.220 ;
        RECT 21.650 118.830 21.820 119.000 ;
        RECT 23.200 118.830 23.370 119.000 ;
        RECT 22.070 118.610 22.950 118.780 ;
        RECT 25.415 119.060 26.295 119.230 ;
        RECT 24.950 118.840 25.120 119.010 ;
        RECT 26.590 118.840 26.760 119.010 ;
        RECT 25.415 118.620 26.295 118.790 ;
        RECT 27.130 118.100 27.390 119.750 ;
        RECT 15.405 116.960 16.285 117.130 ;
        RECT 14.940 116.740 15.110 116.910 ;
        RECT 16.580 116.740 16.750 116.910 ;
        RECT 15.405 116.520 16.285 116.690 ;
        RECT 18.750 116.950 19.630 117.120 ;
        RECT 18.330 116.730 18.500 116.900 ;
        RECT 19.880 116.730 20.050 116.900 ;
        RECT 18.750 116.510 19.630 116.680 ;
        RECT 20.430 115.970 20.690 117.620 ;
        RECT 22.070 116.950 22.950 117.120 ;
        RECT 21.650 116.730 21.820 116.900 ;
        RECT 23.200 116.730 23.370 116.900 ;
        RECT 22.070 116.510 22.950 116.680 ;
        RECT 25.415 116.960 26.295 117.130 ;
        RECT 24.950 116.740 25.120 116.910 ;
        RECT 26.590 116.740 26.760 116.910 ;
        RECT 25.415 116.520 26.295 116.690 ;
        RECT 27.130 116.000 27.390 117.650 ;
        RECT 15.405 114.860 16.285 115.030 ;
        RECT 14.940 114.640 15.110 114.810 ;
        RECT 16.580 114.640 16.750 114.810 ;
        RECT 15.405 114.420 16.285 114.590 ;
        RECT 18.750 114.850 19.630 115.020 ;
        RECT 18.330 114.630 18.500 114.800 ;
        RECT 19.880 114.630 20.050 114.800 ;
        RECT 18.750 114.410 19.630 114.580 ;
        RECT 20.430 113.870 20.690 115.520 ;
        RECT 22.070 114.850 22.950 115.020 ;
        RECT 21.650 114.630 21.820 114.800 ;
        RECT 23.200 114.630 23.370 114.800 ;
        RECT 22.070 114.410 22.950 114.580 ;
        RECT 25.415 114.860 26.295 115.030 ;
        RECT 24.950 114.640 25.120 114.810 ;
        RECT 26.590 114.640 26.760 114.810 ;
        RECT 25.415 114.420 26.295 114.590 ;
        RECT 27.130 113.900 27.390 115.550 ;
        RECT 15.405 112.760 16.285 112.930 ;
        RECT 14.940 112.540 15.110 112.710 ;
        RECT 16.580 112.540 16.750 112.710 ;
        RECT 15.405 112.320 16.285 112.490 ;
        RECT 18.750 112.750 19.630 112.920 ;
        RECT 18.330 112.530 18.500 112.700 ;
        RECT 19.880 112.530 20.050 112.700 ;
        RECT 18.750 112.310 19.630 112.480 ;
        RECT 20.430 111.770 20.690 113.420 ;
        RECT 22.070 112.750 22.950 112.920 ;
        RECT 21.650 112.530 21.820 112.700 ;
        RECT 23.200 112.530 23.370 112.700 ;
        RECT 22.070 112.310 22.950 112.480 ;
        RECT 25.415 112.760 26.295 112.930 ;
        RECT 24.950 112.540 25.120 112.710 ;
        RECT 26.590 112.540 26.760 112.710 ;
        RECT 25.415 112.320 26.295 112.490 ;
        RECT 27.130 111.800 27.390 113.450 ;
        RECT 15.405 110.660 16.285 110.830 ;
        RECT 14.940 110.440 15.110 110.610 ;
        RECT 16.580 110.440 16.750 110.610 ;
        RECT 15.405 110.220 16.285 110.390 ;
        RECT 18.750 110.650 19.630 110.820 ;
        RECT 18.330 110.430 18.500 110.600 ;
        RECT 19.880 110.430 20.050 110.600 ;
        RECT 18.750 110.210 19.630 110.380 ;
        RECT 20.430 109.670 20.690 111.320 ;
        RECT 22.070 110.650 22.950 110.820 ;
        RECT 21.650 110.430 21.820 110.600 ;
        RECT 23.200 110.430 23.370 110.600 ;
        RECT 22.070 110.210 22.950 110.380 ;
        RECT 25.415 110.660 26.295 110.830 ;
        RECT 24.950 110.440 25.120 110.610 ;
        RECT 26.590 110.440 26.760 110.610 ;
        RECT 25.415 110.220 26.295 110.390 ;
        RECT 27.130 109.700 27.390 111.350 ;
        RECT 15.405 108.560 16.285 108.730 ;
        RECT 14.940 108.340 15.110 108.510 ;
        RECT 16.580 108.340 16.750 108.510 ;
        RECT 15.405 108.120 16.285 108.290 ;
        RECT 18.750 108.550 19.630 108.720 ;
        RECT 18.330 108.330 18.500 108.500 ;
        RECT 19.880 108.330 20.050 108.500 ;
        RECT 18.750 108.110 19.630 108.280 ;
        RECT 20.430 107.570 20.690 109.220 ;
        RECT 22.070 108.550 22.950 108.720 ;
        RECT 21.650 108.330 21.820 108.500 ;
        RECT 23.200 108.330 23.370 108.500 ;
        RECT 22.070 108.110 22.950 108.280 ;
        RECT 25.415 108.560 26.295 108.730 ;
        RECT 24.950 108.340 25.120 108.510 ;
        RECT 26.590 108.340 26.760 108.510 ;
        RECT 25.415 108.120 26.295 108.290 ;
        RECT 27.130 107.600 27.390 109.250 ;
        RECT 15.405 106.460 16.285 106.630 ;
        RECT 14.940 106.240 15.110 106.410 ;
        RECT 16.580 106.240 16.750 106.410 ;
        RECT 15.405 106.020 16.285 106.190 ;
        RECT 18.750 106.450 19.630 106.620 ;
        RECT 18.330 106.230 18.500 106.400 ;
        RECT 19.880 106.230 20.050 106.400 ;
        RECT 18.750 106.010 19.630 106.180 ;
        RECT 20.430 105.470 20.690 107.120 ;
        RECT 22.070 106.450 22.950 106.620 ;
        RECT 21.650 106.230 21.820 106.400 ;
        RECT 23.200 106.230 23.370 106.400 ;
        RECT 22.070 106.010 22.950 106.180 ;
        RECT 25.415 106.460 26.295 106.630 ;
        RECT 24.950 106.240 25.120 106.410 ;
        RECT 26.590 106.240 26.760 106.410 ;
        RECT 25.415 106.020 26.295 106.190 ;
        RECT 27.130 105.500 27.390 107.150 ;
        RECT 15.405 104.360 16.285 104.530 ;
        RECT 14.940 104.140 15.110 104.310 ;
        RECT 16.580 104.140 16.750 104.310 ;
        RECT 15.405 103.920 16.285 104.090 ;
        RECT 18.750 104.350 19.630 104.520 ;
        RECT 18.330 104.130 18.500 104.300 ;
        RECT 19.880 104.130 20.050 104.300 ;
        RECT 18.750 103.910 19.630 104.080 ;
        RECT 20.430 103.370 20.690 105.020 ;
        RECT 22.070 104.350 22.950 104.520 ;
        RECT 21.650 104.130 21.820 104.300 ;
        RECT 23.200 104.130 23.370 104.300 ;
        RECT 22.070 103.910 22.950 104.080 ;
        RECT 25.415 104.360 26.295 104.530 ;
        RECT 24.950 104.140 25.120 104.310 ;
        RECT 26.590 104.140 26.760 104.310 ;
        RECT 25.415 103.920 26.295 104.090 ;
        RECT 27.130 103.400 27.390 105.050 ;
        RECT 15.405 102.260 16.285 102.430 ;
        RECT 14.940 102.040 15.110 102.210 ;
        RECT 16.580 102.040 16.750 102.210 ;
        RECT 15.405 101.820 16.285 101.990 ;
        RECT 18.750 102.250 19.630 102.420 ;
        RECT 18.330 102.030 18.500 102.200 ;
        RECT 19.880 102.030 20.050 102.200 ;
        RECT 18.750 101.810 19.630 101.980 ;
        RECT 20.430 101.270 20.690 102.920 ;
        RECT 22.070 102.250 22.950 102.420 ;
        RECT 21.650 102.030 21.820 102.200 ;
        RECT 23.200 102.030 23.370 102.200 ;
        RECT 22.070 101.810 22.950 101.980 ;
        RECT 25.415 102.260 26.295 102.430 ;
        RECT 24.950 102.040 25.120 102.210 ;
        RECT 26.590 102.040 26.760 102.210 ;
        RECT 25.415 101.820 26.295 101.990 ;
        RECT 27.130 101.300 27.390 102.950 ;
        RECT 15.405 100.160 16.285 100.330 ;
        RECT 14.940 99.940 15.110 100.110 ;
        RECT 16.580 99.940 16.750 100.110 ;
        RECT 15.405 99.720 16.285 99.890 ;
        RECT 18.750 100.150 19.630 100.320 ;
        RECT 18.330 99.930 18.500 100.100 ;
        RECT 19.880 99.930 20.050 100.100 ;
        RECT 18.750 99.710 19.630 99.880 ;
        RECT 20.430 99.170 20.690 100.820 ;
        RECT 22.070 100.150 22.950 100.320 ;
        RECT 21.650 99.930 21.820 100.100 ;
        RECT 23.200 99.930 23.370 100.100 ;
        RECT 22.070 99.710 22.950 99.880 ;
        RECT 25.415 100.160 26.295 100.330 ;
        RECT 24.950 99.940 25.120 100.110 ;
        RECT 26.590 99.940 26.760 100.110 ;
        RECT 25.415 99.720 26.295 99.890 ;
        RECT 27.130 99.200 27.390 100.850 ;
        RECT 15.405 98.060 16.285 98.230 ;
        RECT 14.940 97.840 15.110 98.010 ;
        RECT 16.580 97.840 16.750 98.010 ;
        RECT 15.405 97.620 16.285 97.790 ;
        RECT 18.750 98.050 19.630 98.220 ;
        RECT 18.330 97.830 18.500 98.000 ;
        RECT 19.880 97.830 20.050 98.000 ;
        RECT 18.750 97.610 19.630 97.780 ;
        RECT 20.430 97.070 20.690 98.720 ;
        RECT 22.070 98.050 22.950 98.220 ;
        RECT 21.650 97.830 21.820 98.000 ;
        RECT 23.200 97.830 23.370 98.000 ;
        RECT 22.070 97.610 22.950 97.780 ;
        RECT 25.415 98.060 26.295 98.230 ;
        RECT 24.950 97.840 25.120 98.010 ;
        RECT 26.590 97.840 26.760 98.010 ;
        RECT 25.415 97.620 26.295 97.790 ;
        RECT 27.130 97.100 27.390 98.750 ;
        RECT 15.405 95.960 16.285 96.130 ;
        RECT 14.940 95.740 15.110 95.910 ;
        RECT 16.580 95.740 16.750 95.910 ;
        RECT 15.405 95.520 16.285 95.690 ;
        RECT 18.750 95.950 19.630 96.120 ;
        RECT 18.330 95.730 18.500 95.900 ;
        RECT 19.880 95.730 20.050 95.900 ;
        RECT 18.750 95.510 19.630 95.680 ;
        RECT 20.430 94.970 20.690 96.620 ;
        RECT 22.070 95.950 22.950 96.120 ;
        RECT 21.650 95.730 21.820 95.900 ;
        RECT 23.200 95.730 23.370 95.900 ;
        RECT 22.070 95.510 22.950 95.680 ;
        RECT 25.415 95.960 26.295 96.130 ;
        RECT 24.950 95.740 25.120 95.910 ;
        RECT 26.590 95.740 26.760 95.910 ;
        RECT 25.415 95.520 26.295 95.690 ;
        RECT 27.130 95.000 27.390 96.650 ;
        RECT 15.405 93.860 16.285 94.030 ;
        RECT 14.940 93.640 15.110 93.810 ;
        RECT 16.580 93.640 16.750 93.810 ;
        RECT 15.405 93.420 16.285 93.590 ;
        RECT 18.750 93.850 19.630 94.020 ;
        RECT 18.330 93.630 18.500 93.800 ;
        RECT 19.880 93.630 20.050 93.800 ;
        RECT 18.750 93.410 19.630 93.580 ;
        RECT 20.430 92.870 20.690 94.520 ;
        RECT 22.070 93.850 22.950 94.020 ;
        RECT 21.650 93.630 21.820 93.800 ;
        RECT 23.200 93.630 23.370 93.800 ;
        RECT 22.070 93.410 22.950 93.580 ;
        RECT 25.415 93.860 26.295 94.030 ;
        RECT 24.950 93.640 25.120 93.810 ;
        RECT 26.590 93.640 26.760 93.810 ;
        RECT 25.415 93.420 26.295 93.590 ;
        RECT 27.130 92.900 27.390 94.550 ;
        RECT 15.405 91.760 16.285 91.930 ;
        RECT 14.940 91.540 15.110 91.710 ;
        RECT 16.580 91.540 16.750 91.710 ;
        RECT 15.405 91.320 16.285 91.490 ;
        RECT 18.750 91.750 19.630 91.920 ;
        RECT 18.330 91.530 18.500 91.700 ;
        RECT 19.880 91.530 20.050 91.700 ;
        RECT 18.750 91.310 19.630 91.480 ;
        RECT 20.430 90.770 20.690 92.420 ;
        RECT 22.070 91.750 22.950 91.920 ;
        RECT 21.650 91.530 21.820 91.700 ;
        RECT 23.200 91.530 23.370 91.700 ;
        RECT 22.070 91.310 22.950 91.480 ;
        RECT 25.415 91.760 26.295 91.930 ;
        RECT 24.950 91.540 25.120 91.710 ;
        RECT 26.590 91.540 26.760 91.710 ;
        RECT 25.415 91.320 26.295 91.490 ;
        RECT 27.130 90.800 27.390 92.450 ;
        RECT 15.405 89.660 16.285 89.830 ;
        RECT 14.940 89.440 15.110 89.610 ;
        RECT 16.580 89.440 16.750 89.610 ;
        RECT 15.405 89.220 16.285 89.390 ;
        RECT 18.750 89.650 19.630 89.820 ;
        RECT 18.330 89.430 18.500 89.600 ;
        RECT 19.880 89.430 20.050 89.600 ;
        RECT 18.750 89.210 19.630 89.380 ;
        RECT 20.430 88.670 20.690 90.320 ;
        RECT 22.070 89.650 22.950 89.820 ;
        RECT 21.650 89.430 21.820 89.600 ;
        RECT 23.200 89.430 23.370 89.600 ;
        RECT 22.070 89.210 22.950 89.380 ;
        RECT 25.415 89.660 26.295 89.830 ;
        RECT 24.950 89.440 25.120 89.610 ;
        RECT 26.590 89.440 26.760 89.610 ;
        RECT 25.415 89.220 26.295 89.390 ;
        RECT 27.130 88.700 27.390 90.350 ;
        RECT 15.405 87.560 16.285 87.730 ;
        RECT 14.940 87.340 15.110 87.510 ;
        RECT 16.580 87.340 16.750 87.510 ;
        RECT 15.405 87.120 16.285 87.290 ;
        RECT 18.750 87.550 19.630 87.720 ;
        RECT 18.330 87.330 18.500 87.500 ;
        RECT 19.880 87.330 20.050 87.500 ;
        RECT 18.750 87.110 19.630 87.280 ;
        RECT 20.430 86.570 20.690 88.220 ;
        RECT 22.070 87.550 22.950 87.720 ;
        RECT 21.650 87.330 21.820 87.500 ;
        RECT 23.200 87.330 23.370 87.500 ;
        RECT 22.070 87.110 22.950 87.280 ;
        RECT 25.415 87.560 26.295 87.730 ;
        RECT 24.950 87.340 25.120 87.510 ;
        RECT 26.590 87.340 26.760 87.510 ;
        RECT 25.415 87.120 26.295 87.290 ;
        RECT 27.130 86.600 27.390 88.250 ;
        RECT 15.405 85.460 16.285 85.630 ;
        RECT 14.940 85.240 15.110 85.410 ;
        RECT 16.580 85.240 16.750 85.410 ;
        RECT 15.405 85.020 16.285 85.190 ;
        RECT 18.750 85.450 19.630 85.620 ;
        RECT 18.330 85.230 18.500 85.400 ;
        RECT 19.880 85.230 20.050 85.400 ;
        RECT 18.750 85.010 19.630 85.180 ;
        RECT 20.430 84.470 20.690 86.120 ;
        RECT 22.070 85.450 22.950 85.620 ;
        RECT 21.650 85.230 21.820 85.400 ;
        RECT 23.200 85.230 23.370 85.400 ;
        RECT 22.070 85.010 22.950 85.180 ;
        RECT 25.415 85.460 26.295 85.630 ;
        RECT 24.950 85.240 25.120 85.410 ;
        RECT 26.590 85.240 26.760 85.410 ;
        RECT 25.415 85.020 26.295 85.190 ;
        RECT 27.130 84.500 27.390 86.150 ;
        RECT 15.405 83.360 16.285 83.530 ;
        RECT 14.940 83.140 15.110 83.310 ;
        RECT 16.580 83.140 16.750 83.310 ;
        RECT 15.405 82.920 16.285 83.090 ;
        RECT 18.750 83.350 19.630 83.520 ;
        RECT 18.330 83.130 18.500 83.300 ;
        RECT 19.880 83.130 20.050 83.300 ;
        RECT 18.750 82.910 19.630 83.080 ;
        RECT 20.430 82.370 20.690 84.020 ;
        RECT 22.070 83.350 22.950 83.520 ;
        RECT 21.650 83.130 21.820 83.300 ;
        RECT 23.200 83.130 23.370 83.300 ;
        RECT 22.070 82.910 22.950 83.080 ;
        RECT 25.415 83.360 26.295 83.530 ;
        RECT 24.950 83.140 25.120 83.310 ;
        RECT 26.590 83.140 26.760 83.310 ;
        RECT 25.415 82.920 26.295 83.090 ;
        RECT 27.130 82.400 27.390 84.050 ;
        RECT 15.405 81.260 16.285 81.430 ;
        RECT 14.940 81.040 15.110 81.210 ;
        RECT 16.580 81.040 16.750 81.210 ;
        RECT 15.405 80.820 16.285 80.990 ;
        RECT 18.750 81.250 19.630 81.420 ;
        RECT 18.330 81.030 18.500 81.200 ;
        RECT 19.880 81.030 20.050 81.200 ;
        RECT 18.750 80.810 19.630 80.980 ;
        RECT 20.430 80.270 20.690 81.920 ;
        RECT 22.070 81.250 22.950 81.420 ;
        RECT 21.650 81.030 21.820 81.200 ;
        RECT 23.200 81.030 23.370 81.200 ;
        RECT 22.070 80.810 22.950 80.980 ;
        RECT 25.415 81.260 26.295 81.430 ;
        RECT 24.950 81.040 25.120 81.210 ;
        RECT 26.590 81.040 26.760 81.210 ;
        RECT 25.415 80.820 26.295 80.990 ;
        RECT 27.130 80.300 27.390 81.950 ;
        RECT 15.405 79.160 16.285 79.330 ;
        RECT 14.940 78.940 15.110 79.110 ;
        RECT 16.580 78.940 16.750 79.110 ;
        RECT 15.405 78.720 16.285 78.890 ;
        RECT 18.750 79.150 19.630 79.320 ;
        RECT 18.330 78.930 18.500 79.100 ;
        RECT 19.880 78.930 20.050 79.100 ;
        RECT 18.750 78.710 19.630 78.880 ;
        RECT 20.430 78.170 20.690 79.820 ;
        RECT 22.070 79.150 22.950 79.320 ;
        RECT 21.650 78.930 21.820 79.100 ;
        RECT 23.200 78.930 23.370 79.100 ;
        RECT 22.070 78.710 22.950 78.880 ;
        RECT 25.415 79.160 26.295 79.330 ;
        RECT 24.950 78.940 25.120 79.110 ;
        RECT 26.590 78.940 26.760 79.110 ;
        RECT 25.415 78.720 26.295 78.890 ;
        RECT 27.130 78.200 27.390 79.850 ;
        RECT 15.405 77.060 16.285 77.230 ;
        RECT 14.940 76.840 15.110 77.010 ;
        RECT 16.580 76.840 16.750 77.010 ;
        RECT 15.405 76.620 16.285 76.790 ;
        RECT 18.750 77.050 19.630 77.220 ;
        RECT 18.330 76.830 18.500 77.000 ;
        RECT 19.880 76.830 20.050 77.000 ;
        RECT 18.750 76.610 19.630 76.780 ;
        RECT 20.430 76.070 20.690 77.720 ;
        RECT 22.070 77.050 22.950 77.220 ;
        RECT 21.650 76.830 21.820 77.000 ;
        RECT 23.200 76.830 23.370 77.000 ;
        RECT 22.070 76.610 22.950 76.780 ;
        RECT 25.415 77.060 26.295 77.230 ;
        RECT 24.950 76.840 25.120 77.010 ;
        RECT 26.590 76.840 26.760 77.010 ;
        RECT 25.415 76.620 26.295 76.790 ;
        RECT 27.130 76.100 27.390 77.750 ;
        RECT 15.405 74.960 16.285 75.130 ;
        RECT 14.940 74.740 15.110 74.910 ;
        RECT 16.580 74.740 16.750 74.910 ;
        RECT 15.405 74.520 16.285 74.690 ;
        RECT 18.750 74.950 19.630 75.120 ;
        RECT 18.330 74.730 18.500 74.900 ;
        RECT 19.880 74.730 20.050 74.900 ;
        RECT 18.750 74.510 19.630 74.680 ;
        RECT 20.430 73.970 20.690 75.620 ;
        RECT 22.070 74.950 22.950 75.120 ;
        RECT 21.650 74.730 21.820 74.900 ;
        RECT 23.200 74.730 23.370 74.900 ;
        RECT 22.070 74.510 22.950 74.680 ;
        RECT 25.415 74.960 26.295 75.130 ;
        RECT 24.950 74.740 25.120 74.910 ;
        RECT 26.590 74.740 26.760 74.910 ;
        RECT 25.415 74.520 26.295 74.690 ;
        RECT 27.130 74.000 27.390 75.650 ;
        RECT 15.405 72.860 16.285 73.030 ;
        RECT 14.940 72.640 15.110 72.810 ;
        RECT 16.580 72.640 16.750 72.810 ;
        RECT 15.405 72.420 16.285 72.590 ;
        RECT 18.750 72.850 19.630 73.020 ;
        RECT 18.330 72.630 18.500 72.800 ;
        RECT 19.880 72.630 20.050 72.800 ;
        RECT 18.750 72.410 19.630 72.580 ;
        RECT 20.430 71.870 20.690 73.520 ;
        RECT 22.070 72.850 22.950 73.020 ;
        RECT 21.650 72.630 21.820 72.800 ;
        RECT 23.200 72.630 23.370 72.800 ;
        RECT 22.070 72.410 22.950 72.580 ;
        RECT 25.415 72.860 26.295 73.030 ;
        RECT 24.950 72.640 25.120 72.810 ;
        RECT 26.590 72.640 26.760 72.810 ;
        RECT 25.415 72.420 26.295 72.590 ;
        RECT 27.130 71.900 27.390 73.550 ;
        RECT 15.405 70.760 16.285 70.930 ;
        RECT 14.940 70.540 15.110 70.710 ;
        RECT 16.580 70.540 16.750 70.710 ;
        RECT 15.405 70.320 16.285 70.490 ;
        RECT 18.750 70.750 19.630 70.920 ;
        RECT 18.330 70.530 18.500 70.700 ;
        RECT 19.880 70.530 20.050 70.700 ;
        RECT 18.750 70.310 19.630 70.480 ;
        RECT 20.430 69.770 20.690 71.420 ;
        RECT 22.070 70.750 22.950 70.920 ;
        RECT 21.650 70.530 21.820 70.700 ;
        RECT 23.200 70.530 23.370 70.700 ;
        RECT 22.070 70.310 22.950 70.480 ;
        RECT 25.415 70.760 26.295 70.930 ;
        RECT 24.950 70.540 25.120 70.710 ;
        RECT 26.590 70.540 26.760 70.710 ;
        RECT 25.415 70.320 26.295 70.490 ;
        RECT 27.130 69.800 27.390 71.450 ;
        RECT 15.405 68.660 16.285 68.830 ;
        RECT 14.940 68.440 15.110 68.610 ;
        RECT 16.580 68.440 16.750 68.610 ;
        RECT 15.405 68.220 16.285 68.390 ;
        RECT 18.750 68.650 19.630 68.820 ;
        RECT 18.330 68.430 18.500 68.600 ;
        RECT 19.880 68.430 20.050 68.600 ;
        RECT 18.750 68.210 19.630 68.380 ;
        RECT 20.430 67.670 20.690 69.320 ;
        RECT 22.070 68.650 22.950 68.820 ;
        RECT 21.650 68.430 21.820 68.600 ;
        RECT 23.200 68.430 23.370 68.600 ;
        RECT 22.070 68.210 22.950 68.380 ;
        RECT 25.415 68.660 26.295 68.830 ;
        RECT 24.950 68.440 25.120 68.610 ;
        RECT 26.590 68.440 26.760 68.610 ;
        RECT 25.415 68.220 26.295 68.390 ;
        RECT 27.130 67.700 27.390 69.350 ;
        RECT 15.405 66.560 16.285 66.730 ;
        RECT 14.940 66.340 15.110 66.510 ;
        RECT 16.580 66.340 16.750 66.510 ;
        RECT 15.405 66.120 16.285 66.290 ;
        RECT 18.750 66.550 19.630 66.720 ;
        RECT 18.330 66.330 18.500 66.500 ;
        RECT 19.880 66.330 20.050 66.500 ;
        RECT 18.750 66.110 19.630 66.280 ;
        RECT 20.430 65.570 20.690 67.220 ;
        RECT 22.070 66.550 22.950 66.720 ;
        RECT 21.650 66.330 21.820 66.500 ;
        RECT 23.200 66.330 23.370 66.500 ;
        RECT 22.070 66.110 22.950 66.280 ;
        RECT 25.415 66.560 26.295 66.730 ;
        RECT 24.950 66.340 25.120 66.510 ;
        RECT 26.590 66.340 26.760 66.510 ;
        RECT 25.415 66.120 26.295 66.290 ;
        RECT 27.130 65.600 27.390 67.250 ;
        RECT 15.405 64.460 16.285 64.630 ;
        RECT 14.940 64.240 15.110 64.410 ;
        RECT 16.580 64.240 16.750 64.410 ;
        RECT 15.405 64.020 16.285 64.190 ;
        RECT 18.750 64.450 19.630 64.620 ;
        RECT 18.330 64.230 18.500 64.400 ;
        RECT 19.880 64.230 20.050 64.400 ;
        RECT 18.750 64.010 19.630 64.180 ;
        RECT 20.430 63.470 20.690 65.120 ;
        RECT 22.070 64.450 22.950 64.620 ;
        RECT 21.650 64.230 21.820 64.400 ;
        RECT 23.200 64.230 23.370 64.400 ;
        RECT 22.070 64.010 22.950 64.180 ;
        RECT 25.415 64.460 26.295 64.630 ;
        RECT 24.950 64.240 25.120 64.410 ;
        RECT 26.590 64.240 26.760 64.410 ;
        RECT 25.415 64.020 26.295 64.190 ;
        RECT 27.130 63.500 27.390 65.150 ;
        RECT 15.405 62.360 16.285 62.530 ;
        RECT 14.940 62.140 15.110 62.310 ;
        RECT 16.580 62.140 16.750 62.310 ;
        RECT 15.405 61.920 16.285 62.090 ;
        RECT 18.750 62.350 19.630 62.520 ;
        RECT 18.330 62.130 18.500 62.300 ;
        RECT 19.880 62.130 20.050 62.300 ;
        RECT 18.750 61.910 19.630 62.080 ;
        RECT 20.430 61.370 20.690 63.020 ;
        RECT 22.070 62.350 22.950 62.520 ;
        RECT 21.650 62.130 21.820 62.300 ;
        RECT 23.200 62.130 23.370 62.300 ;
        RECT 22.070 61.910 22.950 62.080 ;
        RECT 25.415 62.360 26.295 62.530 ;
        RECT 24.950 62.140 25.120 62.310 ;
        RECT 26.590 62.140 26.760 62.310 ;
        RECT 25.415 61.920 26.295 62.090 ;
        RECT 27.130 61.400 27.390 63.050 ;
        RECT 15.405 60.260 16.285 60.430 ;
        RECT 14.940 60.040 15.110 60.210 ;
        RECT 16.580 60.040 16.750 60.210 ;
        RECT 15.405 59.820 16.285 59.990 ;
        RECT 18.750 60.250 19.630 60.420 ;
        RECT 18.330 60.030 18.500 60.200 ;
        RECT 19.880 60.030 20.050 60.200 ;
        RECT 18.750 59.810 19.630 59.980 ;
        RECT 20.430 59.270 20.690 60.920 ;
        RECT 22.070 60.250 22.950 60.420 ;
        RECT 21.650 60.030 21.820 60.200 ;
        RECT 23.200 60.030 23.370 60.200 ;
        RECT 22.070 59.810 22.950 59.980 ;
        RECT 25.415 60.260 26.295 60.430 ;
        RECT 24.950 60.040 25.120 60.210 ;
        RECT 26.590 60.040 26.760 60.210 ;
        RECT 25.415 59.820 26.295 59.990 ;
        RECT 27.130 59.300 27.390 60.950 ;
        RECT 15.405 58.160 16.285 58.330 ;
        RECT 14.940 57.940 15.110 58.110 ;
        RECT 16.580 57.940 16.750 58.110 ;
        RECT 15.405 57.720 16.285 57.890 ;
        RECT 18.750 58.150 19.630 58.320 ;
        RECT 18.330 57.930 18.500 58.100 ;
        RECT 19.880 57.930 20.050 58.100 ;
        RECT 18.750 57.710 19.630 57.880 ;
        RECT 20.430 57.170 20.690 58.820 ;
        RECT 22.070 58.150 22.950 58.320 ;
        RECT 21.650 57.930 21.820 58.100 ;
        RECT 23.200 57.930 23.370 58.100 ;
        RECT 22.070 57.710 22.950 57.880 ;
        RECT 25.415 58.160 26.295 58.330 ;
        RECT 24.950 57.940 25.120 58.110 ;
        RECT 26.590 57.940 26.760 58.110 ;
        RECT 25.415 57.720 26.295 57.890 ;
        RECT 27.130 57.200 27.390 58.850 ;
        RECT 15.405 56.060 16.285 56.230 ;
        RECT 14.940 55.840 15.110 56.010 ;
        RECT 16.580 55.840 16.750 56.010 ;
        RECT 15.405 55.620 16.285 55.790 ;
        RECT 18.750 56.050 19.630 56.220 ;
        RECT 18.330 55.830 18.500 56.000 ;
        RECT 19.880 55.830 20.050 56.000 ;
        RECT 18.750 55.610 19.630 55.780 ;
        RECT 20.430 55.070 20.690 56.720 ;
        RECT 22.070 56.050 22.950 56.220 ;
        RECT 21.650 55.830 21.820 56.000 ;
        RECT 23.200 55.830 23.370 56.000 ;
        RECT 22.070 55.610 22.950 55.780 ;
        RECT 25.415 56.060 26.295 56.230 ;
        RECT 24.950 55.840 25.120 56.010 ;
        RECT 26.590 55.840 26.760 56.010 ;
        RECT 25.415 55.620 26.295 55.790 ;
        RECT 27.130 55.100 27.390 56.750 ;
        RECT 15.405 53.960 16.285 54.130 ;
        RECT 14.940 53.740 15.110 53.910 ;
        RECT 16.580 53.740 16.750 53.910 ;
        RECT 15.405 53.520 16.285 53.690 ;
        RECT 18.750 53.950 19.630 54.120 ;
        RECT 18.330 53.730 18.500 53.900 ;
        RECT 19.880 53.730 20.050 53.900 ;
        RECT 18.750 53.510 19.630 53.680 ;
        RECT 20.430 52.970 20.690 54.620 ;
        RECT 22.070 53.950 22.950 54.120 ;
        RECT 21.650 53.730 21.820 53.900 ;
        RECT 23.200 53.730 23.370 53.900 ;
        RECT 22.070 53.510 22.950 53.680 ;
        RECT 25.415 53.960 26.295 54.130 ;
        RECT 24.950 53.740 25.120 53.910 ;
        RECT 26.590 53.740 26.760 53.910 ;
        RECT 25.415 53.520 26.295 53.690 ;
        RECT 27.130 53.000 27.390 54.650 ;
        RECT 15.405 51.860 16.285 52.030 ;
        RECT 14.940 51.640 15.110 51.810 ;
        RECT 16.580 51.640 16.750 51.810 ;
        RECT 15.405 51.420 16.285 51.590 ;
        RECT 18.750 51.850 19.630 52.020 ;
        RECT 18.330 51.630 18.500 51.800 ;
        RECT 19.880 51.630 20.050 51.800 ;
        RECT 18.750 51.410 19.630 51.580 ;
        RECT 20.430 50.870 20.690 52.520 ;
        RECT 22.070 51.850 22.950 52.020 ;
        RECT 21.650 51.630 21.820 51.800 ;
        RECT 23.200 51.630 23.370 51.800 ;
        RECT 22.070 51.410 22.950 51.580 ;
        RECT 25.415 51.860 26.295 52.030 ;
        RECT 24.950 51.640 25.120 51.810 ;
        RECT 26.590 51.640 26.760 51.810 ;
        RECT 25.415 51.420 26.295 51.590 ;
        RECT 27.130 50.900 27.390 52.550 ;
        RECT 15.405 49.760 16.285 49.930 ;
        RECT 14.940 49.540 15.110 49.710 ;
        RECT 16.580 49.540 16.750 49.710 ;
        RECT 15.405 49.320 16.285 49.490 ;
        RECT 18.750 49.750 19.630 49.920 ;
        RECT 18.330 49.530 18.500 49.700 ;
        RECT 19.880 49.530 20.050 49.700 ;
        RECT 18.750 49.310 19.630 49.480 ;
        RECT 20.430 48.770 20.690 50.420 ;
        RECT 22.070 49.750 22.950 49.920 ;
        RECT 21.650 49.530 21.820 49.700 ;
        RECT 23.200 49.530 23.370 49.700 ;
        RECT 22.070 49.310 22.950 49.480 ;
        RECT 25.415 49.760 26.295 49.930 ;
        RECT 24.950 49.540 25.120 49.710 ;
        RECT 26.590 49.540 26.760 49.710 ;
        RECT 25.415 49.320 26.295 49.490 ;
        RECT 27.130 48.800 27.390 50.450 ;
        RECT 15.405 47.660 16.285 47.830 ;
        RECT 14.940 47.440 15.110 47.610 ;
        RECT 16.580 47.440 16.750 47.610 ;
        RECT 15.405 47.220 16.285 47.390 ;
        RECT 18.750 47.650 19.630 47.820 ;
        RECT 18.330 47.430 18.500 47.600 ;
        RECT 19.880 47.430 20.050 47.600 ;
        RECT 18.750 47.210 19.630 47.380 ;
        RECT 20.430 46.670 20.690 48.320 ;
        RECT 22.070 47.650 22.950 47.820 ;
        RECT 21.650 47.430 21.820 47.600 ;
        RECT 23.200 47.430 23.370 47.600 ;
        RECT 22.070 47.210 22.950 47.380 ;
        RECT 25.415 47.660 26.295 47.830 ;
        RECT 24.950 47.440 25.120 47.610 ;
        RECT 26.590 47.440 26.760 47.610 ;
        RECT 25.415 47.220 26.295 47.390 ;
        RECT 27.130 46.700 27.390 48.350 ;
        RECT 15.405 45.560 16.285 45.730 ;
        RECT 14.940 45.340 15.110 45.510 ;
        RECT 16.580 45.340 16.750 45.510 ;
        RECT 15.405 45.120 16.285 45.290 ;
        RECT 18.750 45.550 19.630 45.720 ;
        RECT 18.330 45.330 18.500 45.500 ;
        RECT 19.880 45.330 20.050 45.500 ;
        RECT 18.750 45.110 19.630 45.280 ;
        RECT 20.430 44.570 20.690 46.220 ;
        RECT 22.070 45.550 22.950 45.720 ;
        RECT 21.650 45.330 21.820 45.500 ;
        RECT 23.200 45.330 23.370 45.500 ;
        RECT 22.070 45.110 22.950 45.280 ;
        RECT 25.415 45.560 26.295 45.730 ;
        RECT 24.950 45.340 25.120 45.510 ;
        RECT 26.590 45.340 26.760 45.510 ;
        RECT 25.415 45.120 26.295 45.290 ;
        RECT 27.130 44.600 27.390 46.250 ;
        RECT 15.405 43.460 16.285 43.630 ;
        RECT 14.940 43.240 15.110 43.410 ;
        RECT 16.580 43.240 16.750 43.410 ;
        RECT 15.405 43.020 16.285 43.190 ;
        RECT 18.750 43.450 19.630 43.620 ;
        RECT 18.330 43.230 18.500 43.400 ;
        RECT 19.880 43.230 20.050 43.400 ;
        RECT 18.750 43.010 19.630 43.180 ;
        RECT 20.430 42.470 20.690 44.120 ;
        RECT 22.070 43.450 22.950 43.620 ;
        RECT 21.650 43.230 21.820 43.400 ;
        RECT 23.200 43.230 23.370 43.400 ;
        RECT 22.070 43.010 22.950 43.180 ;
        RECT 25.415 43.460 26.295 43.630 ;
        RECT 24.950 43.240 25.120 43.410 ;
        RECT 26.590 43.240 26.760 43.410 ;
        RECT 25.415 43.020 26.295 43.190 ;
        RECT 27.130 42.500 27.390 44.150 ;
        RECT 15.405 41.360 16.285 41.530 ;
        RECT 14.940 41.140 15.110 41.310 ;
        RECT 16.580 41.140 16.750 41.310 ;
        RECT 15.405 40.920 16.285 41.090 ;
        RECT 18.750 41.350 19.630 41.520 ;
        RECT 18.330 41.130 18.500 41.300 ;
        RECT 19.880 41.130 20.050 41.300 ;
        RECT 18.750 40.910 19.630 41.080 ;
        RECT 20.430 40.370 20.690 42.020 ;
        RECT 22.070 41.350 22.950 41.520 ;
        RECT 21.650 41.130 21.820 41.300 ;
        RECT 23.200 41.130 23.370 41.300 ;
        RECT 22.070 40.910 22.950 41.080 ;
        RECT 25.415 41.360 26.295 41.530 ;
        RECT 24.950 41.140 25.120 41.310 ;
        RECT 26.590 41.140 26.760 41.310 ;
        RECT 25.415 40.920 26.295 41.090 ;
        RECT 27.130 40.400 27.390 42.050 ;
        RECT 15.405 39.260 16.285 39.430 ;
        RECT 14.940 39.040 15.110 39.210 ;
        RECT 16.580 39.040 16.750 39.210 ;
        RECT 15.405 38.820 16.285 38.990 ;
        RECT 18.750 39.250 19.630 39.420 ;
        RECT 18.330 39.030 18.500 39.200 ;
        RECT 19.880 39.030 20.050 39.200 ;
        RECT 18.750 38.810 19.630 38.980 ;
        RECT 20.430 38.270 20.690 39.920 ;
        RECT 22.070 39.250 22.950 39.420 ;
        RECT 21.650 39.030 21.820 39.200 ;
        RECT 23.200 39.030 23.370 39.200 ;
        RECT 22.070 38.810 22.950 38.980 ;
        RECT 25.415 39.260 26.295 39.430 ;
        RECT 24.950 39.040 25.120 39.210 ;
        RECT 26.590 39.040 26.760 39.210 ;
        RECT 25.415 38.820 26.295 38.990 ;
        RECT 27.130 38.300 27.390 39.950 ;
        RECT 15.405 37.160 16.285 37.330 ;
        RECT 14.940 36.940 15.110 37.110 ;
        RECT 16.580 36.940 16.750 37.110 ;
        RECT 15.405 36.720 16.285 36.890 ;
        RECT 18.750 37.150 19.630 37.320 ;
        RECT 18.330 36.930 18.500 37.100 ;
        RECT 19.880 36.930 20.050 37.100 ;
        RECT 18.750 36.710 19.630 36.880 ;
        RECT 20.430 36.170 20.690 37.820 ;
        RECT 22.070 37.150 22.950 37.320 ;
        RECT 21.650 36.930 21.820 37.100 ;
        RECT 23.200 36.930 23.370 37.100 ;
        RECT 22.070 36.710 22.950 36.880 ;
        RECT 25.415 37.160 26.295 37.330 ;
        RECT 24.950 36.940 25.120 37.110 ;
        RECT 26.590 36.940 26.760 37.110 ;
        RECT 25.415 36.720 26.295 36.890 ;
        RECT 27.130 36.200 27.390 37.850 ;
        RECT 15.405 35.060 16.285 35.230 ;
        RECT 14.940 34.840 15.110 35.010 ;
        RECT 16.580 34.840 16.750 35.010 ;
        RECT 15.405 34.620 16.285 34.790 ;
        RECT 18.750 35.050 19.630 35.220 ;
        RECT 18.330 34.830 18.500 35.000 ;
        RECT 19.880 34.830 20.050 35.000 ;
        RECT 18.750 34.610 19.630 34.780 ;
        RECT 20.430 34.070 20.690 35.720 ;
        RECT 22.070 35.050 22.950 35.220 ;
        RECT 21.650 34.830 21.820 35.000 ;
        RECT 23.200 34.830 23.370 35.000 ;
        RECT 22.070 34.610 22.950 34.780 ;
        RECT 25.415 35.060 26.295 35.230 ;
        RECT 24.950 34.840 25.120 35.010 ;
        RECT 26.590 34.840 26.760 35.010 ;
        RECT 25.415 34.620 26.295 34.790 ;
        RECT 27.130 34.100 27.390 35.750 ;
        RECT 15.405 32.960 16.285 33.130 ;
        RECT 14.940 32.740 15.110 32.910 ;
        RECT 16.580 32.740 16.750 32.910 ;
        RECT 15.405 32.520 16.285 32.690 ;
        RECT 18.750 32.950 19.630 33.120 ;
        RECT 18.330 32.730 18.500 32.900 ;
        RECT 19.880 32.730 20.050 32.900 ;
        RECT 18.750 32.510 19.630 32.680 ;
        RECT 20.430 31.970 20.690 33.620 ;
        RECT 22.070 32.950 22.950 33.120 ;
        RECT 21.650 32.730 21.820 32.900 ;
        RECT 23.200 32.730 23.370 32.900 ;
        RECT 22.070 32.510 22.950 32.680 ;
        RECT 25.415 32.960 26.295 33.130 ;
        RECT 24.950 32.740 25.120 32.910 ;
        RECT 26.590 32.740 26.760 32.910 ;
        RECT 25.415 32.520 26.295 32.690 ;
        RECT 27.130 32.000 27.390 33.650 ;
        RECT 15.405 30.860 16.285 31.030 ;
        RECT 14.940 30.640 15.110 30.810 ;
        RECT 16.580 30.640 16.750 30.810 ;
        RECT 15.405 30.420 16.285 30.590 ;
        RECT 18.750 30.850 19.630 31.020 ;
        RECT 18.330 30.630 18.500 30.800 ;
        RECT 19.880 30.630 20.050 30.800 ;
        RECT 18.750 30.410 19.630 30.580 ;
        RECT 20.430 29.870 20.690 31.520 ;
        RECT 22.070 30.850 22.950 31.020 ;
        RECT 21.650 30.630 21.820 30.800 ;
        RECT 23.200 30.630 23.370 30.800 ;
        RECT 22.070 30.410 22.950 30.580 ;
        RECT 25.415 30.860 26.295 31.030 ;
        RECT 24.950 30.640 25.120 30.810 ;
        RECT 26.590 30.640 26.760 30.810 ;
        RECT 25.415 30.420 26.295 30.590 ;
        RECT 27.130 29.900 27.390 31.550 ;
        RECT 15.405 28.760 16.285 28.930 ;
        RECT 14.940 28.540 15.110 28.710 ;
        RECT 16.580 28.540 16.750 28.710 ;
        RECT 15.405 28.320 16.285 28.490 ;
        RECT 18.750 28.750 19.630 28.920 ;
        RECT 18.330 28.530 18.500 28.700 ;
        RECT 19.880 28.530 20.050 28.700 ;
        RECT 18.750 28.310 19.630 28.480 ;
        RECT 20.430 27.770 20.690 29.420 ;
        RECT 22.070 28.750 22.950 28.920 ;
        RECT 21.650 28.530 21.820 28.700 ;
        RECT 23.200 28.530 23.370 28.700 ;
        RECT 22.070 28.310 22.950 28.480 ;
        RECT 25.415 28.760 26.295 28.930 ;
        RECT 24.950 28.540 25.120 28.710 ;
        RECT 26.590 28.540 26.760 28.710 ;
        RECT 25.415 28.320 26.295 28.490 ;
        RECT 27.130 27.800 27.390 29.450 ;
        RECT 15.405 26.660 16.285 26.830 ;
        RECT 14.940 26.440 15.110 26.610 ;
        RECT 16.580 26.440 16.750 26.610 ;
        RECT 15.405 26.220 16.285 26.390 ;
        RECT 18.750 26.650 19.630 26.820 ;
        RECT 18.330 26.430 18.500 26.600 ;
        RECT 19.880 26.430 20.050 26.600 ;
        RECT 18.750 26.210 19.630 26.380 ;
        RECT 20.430 25.670 20.690 27.320 ;
        RECT 22.070 26.650 22.950 26.820 ;
        RECT 21.650 26.430 21.820 26.600 ;
        RECT 23.200 26.430 23.370 26.600 ;
        RECT 22.070 26.210 22.950 26.380 ;
        RECT 25.415 26.660 26.295 26.830 ;
        RECT 24.950 26.440 25.120 26.610 ;
        RECT 26.590 26.440 26.760 26.610 ;
        RECT 25.415 26.220 26.295 26.390 ;
        RECT 27.130 25.700 27.390 27.350 ;
        RECT 15.405 24.560 16.285 24.730 ;
        RECT 14.940 24.340 15.110 24.510 ;
        RECT 16.580 24.340 16.750 24.510 ;
        RECT 15.405 24.120 16.285 24.290 ;
        RECT 18.750 24.550 19.630 24.720 ;
        RECT 18.330 24.330 18.500 24.500 ;
        RECT 19.880 24.330 20.050 24.500 ;
        RECT 18.750 24.110 19.630 24.280 ;
        RECT 20.430 23.570 20.690 25.220 ;
        RECT 22.070 24.550 22.950 24.720 ;
        RECT 21.650 24.330 21.820 24.500 ;
        RECT 23.200 24.330 23.370 24.500 ;
        RECT 22.070 24.110 22.950 24.280 ;
        RECT 25.415 24.560 26.295 24.730 ;
        RECT 24.950 24.340 25.120 24.510 ;
        RECT 26.590 24.340 26.760 24.510 ;
        RECT 25.415 24.120 26.295 24.290 ;
        RECT 27.130 23.600 27.390 25.250 ;
        RECT 15.405 22.460 16.285 22.630 ;
        RECT 14.940 22.240 15.110 22.410 ;
        RECT 16.580 22.240 16.750 22.410 ;
        RECT 15.405 22.020 16.285 22.190 ;
        RECT 18.750 22.450 19.630 22.620 ;
        RECT 18.330 22.230 18.500 22.400 ;
        RECT 19.880 22.230 20.050 22.400 ;
        RECT 18.750 22.010 19.630 22.180 ;
        RECT 20.430 21.470 20.690 23.120 ;
        RECT 22.070 22.450 22.950 22.620 ;
        RECT 21.650 22.230 21.820 22.400 ;
        RECT 23.200 22.230 23.370 22.400 ;
        RECT 22.070 22.010 22.950 22.180 ;
        RECT 25.415 22.460 26.295 22.630 ;
        RECT 24.950 22.240 25.120 22.410 ;
        RECT 26.590 22.240 26.760 22.410 ;
        RECT 25.415 22.020 26.295 22.190 ;
        RECT 27.130 21.500 27.390 23.150 ;
        RECT 15.405 20.360 16.285 20.530 ;
        RECT 14.940 20.140 15.110 20.310 ;
        RECT 16.580 20.140 16.750 20.310 ;
        RECT 15.405 19.920 16.285 20.090 ;
        RECT 18.750 20.350 19.630 20.520 ;
        RECT 18.330 20.130 18.500 20.300 ;
        RECT 19.880 20.130 20.050 20.300 ;
        RECT 18.750 19.910 19.630 20.080 ;
        RECT 20.430 19.370 20.690 21.020 ;
        RECT 22.070 20.350 22.950 20.520 ;
        RECT 21.650 20.130 21.820 20.300 ;
        RECT 23.200 20.130 23.370 20.300 ;
        RECT 22.070 19.910 22.950 20.080 ;
        RECT 25.415 20.360 26.295 20.530 ;
        RECT 24.950 20.140 25.120 20.310 ;
        RECT 26.590 20.140 26.760 20.310 ;
        RECT 25.415 19.920 26.295 20.090 ;
        RECT 27.130 19.400 27.390 21.050 ;
        RECT 15.405 18.260 16.285 18.430 ;
        RECT 14.940 18.040 15.110 18.210 ;
        RECT 16.580 18.040 16.750 18.210 ;
        RECT 15.405 17.820 16.285 17.990 ;
        RECT 18.750 18.250 19.630 18.420 ;
        RECT 18.330 18.030 18.500 18.200 ;
        RECT 19.880 18.030 20.050 18.200 ;
        RECT 18.750 17.810 19.630 17.980 ;
        RECT 20.430 17.270 20.690 18.920 ;
        RECT 22.070 18.250 22.950 18.420 ;
        RECT 21.650 18.030 21.820 18.200 ;
        RECT 23.200 18.030 23.370 18.200 ;
        RECT 22.070 17.810 22.950 17.980 ;
        RECT 25.415 18.260 26.295 18.430 ;
        RECT 24.950 18.040 25.120 18.210 ;
        RECT 26.590 18.040 26.760 18.210 ;
        RECT 25.415 17.820 26.295 17.990 ;
        RECT 27.130 17.300 27.390 18.950 ;
        RECT 15.405 16.160 16.285 16.330 ;
        RECT 14.940 15.940 15.110 16.110 ;
        RECT 16.580 15.940 16.750 16.110 ;
        RECT 15.405 15.720 16.285 15.890 ;
        RECT 18.750 16.150 19.630 16.320 ;
        RECT 18.330 15.930 18.500 16.100 ;
        RECT 19.880 15.930 20.050 16.100 ;
        RECT 18.750 15.710 19.630 15.880 ;
        RECT 20.430 15.170 20.690 16.820 ;
        RECT 22.070 16.150 22.950 16.320 ;
        RECT 21.650 15.930 21.820 16.100 ;
        RECT 23.200 15.930 23.370 16.100 ;
        RECT 22.070 15.710 22.950 15.880 ;
        RECT 25.415 16.160 26.295 16.330 ;
        RECT 24.950 15.940 25.120 16.110 ;
        RECT 26.590 15.940 26.760 16.110 ;
        RECT 25.415 15.720 26.295 15.890 ;
        RECT 27.130 15.200 27.390 16.850 ;
        RECT 15.405 14.060 16.285 14.230 ;
        RECT 14.940 13.840 15.110 14.010 ;
        RECT 16.580 13.840 16.750 14.010 ;
        RECT 15.405 13.620 16.285 13.790 ;
        RECT 18.750 14.050 19.630 14.220 ;
        RECT 18.330 13.830 18.500 14.000 ;
        RECT 19.880 13.830 20.050 14.000 ;
        RECT 18.750 13.610 19.630 13.780 ;
        RECT 20.430 13.070 20.690 14.720 ;
        RECT 22.070 14.050 22.950 14.220 ;
        RECT 21.650 13.830 21.820 14.000 ;
        RECT 23.200 13.830 23.370 14.000 ;
        RECT 22.070 13.610 22.950 13.780 ;
        RECT 25.415 14.060 26.295 14.230 ;
        RECT 24.950 13.840 25.120 14.010 ;
        RECT 26.590 13.840 26.760 14.010 ;
        RECT 25.415 13.620 26.295 13.790 ;
        RECT 27.130 13.100 27.390 14.750 ;
        RECT 15.405 11.960 16.285 12.130 ;
        RECT 14.940 11.740 15.110 11.910 ;
        RECT 16.580 11.740 16.750 11.910 ;
        RECT 15.405 11.520 16.285 11.690 ;
        RECT 18.750 11.950 19.630 12.120 ;
        RECT 18.330 11.730 18.500 11.900 ;
        RECT 19.880 11.730 20.050 11.900 ;
        RECT 18.750 11.510 19.630 11.680 ;
        RECT 20.430 10.970 20.690 12.620 ;
        RECT 22.070 11.950 22.950 12.120 ;
        RECT 21.650 11.730 21.820 11.900 ;
        RECT 23.200 11.730 23.370 11.900 ;
        RECT 22.070 11.510 22.950 11.680 ;
        RECT 25.415 11.960 26.295 12.130 ;
        RECT 24.950 11.740 25.120 11.910 ;
        RECT 26.590 11.740 26.760 11.910 ;
        RECT 25.415 11.520 26.295 11.690 ;
        RECT 27.130 11.000 27.390 12.650 ;
      LAYER met1 ;
        RECT 20.950 220.760 21.320 220.770 ;
        RECT 14.250 220.600 14.600 220.710 ;
        RECT 14.250 220.330 16.370 220.600 ;
        RECT 14.250 218.500 14.600 220.330 ;
        RECT 14.850 219.500 15.170 219.830 ;
        RECT 15.330 219.800 16.360 220.330 ;
        RECT 17.090 219.830 17.820 220.700 ;
        RECT 20.380 220.590 21.320 220.760 ;
        RECT 20.380 220.530 23.010 220.590 ;
        RECT 18.690 220.320 23.010 220.530 ;
        RECT 18.690 220.260 21.320 220.320 ;
        RECT 15.345 219.770 16.345 219.800 ;
        RECT 15.345 219.540 16.345 219.560 ;
        RECT 15.330 219.240 16.370 219.540 ;
        RECT 16.520 219.500 18.550 219.830 ;
        RECT 18.690 219.710 19.690 220.260 ;
        RECT 19.870 219.800 20.130 219.830 ;
        RECT 18.690 219.540 19.690 219.550 ;
        RECT 18.690 219.330 19.700 219.540 ;
        RECT 19.850 219.510 20.130 219.800 ;
        RECT 19.870 219.490 20.130 219.510 ;
        RECT 18.550 219.240 19.700 219.330 ;
        RECT 15.330 219.100 19.700 219.240 ;
        RECT 16.320 219.080 19.700 219.100 ;
        RECT 14.250 218.230 16.370 218.500 ;
        RECT 14.250 216.400 14.600 218.230 ;
        RECT 14.850 217.400 15.170 217.730 ;
        RECT 15.330 217.700 16.360 218.230 ;
        RECT 17.090 217.730 17.820 219.080 ;
        RECT 20.380 218.490 21.320 220.260 ;
        RECT 21.570 219.860 21.830 219.890 ;
        RECT 21.570 219.570 21.850 219.860 ;
        RECT 22.010 219.770 23.010 220.320 ;
        RECT 23.880 219.890 24.610 220.760 ;
        RECT 27.100 220.660 27.450 220.770 ;
        RECT 25.330 220.390 27.450 220.660 ;
        RECT 22.010 219.600 23.010 219.610 ;
        RECT 21.570 219.550 21.830 219.570 ;
        RECT 22.000 219.390 23.010 219.600 ;
        RECT 23.150 219.560 25.180 219.890 ;
        RECT 25.340 219.860 26.370 220.390 ;
        RECT 25.355 219.830 26.355 219.860 ;
        RECT 25.355 219.600 26.355 219.620 ;
        RECT 22.000 219.300 23.150 219.390 ;
        RECT 25.330 219.300 26.370 219.600 ;
        RECT 26.530 219.560 26.850 219.890 ;
        RECT 22.000 219.160 26.370 219.300 ;
        RECT 22.000 219.140 25.380 219.160 ;
        RECT 20.380 218.430 23.010 218.490 ;
        RECT 18.690 218.220 23.010 218.430 ;
        RECT 18.690 218.160 21.320 218.220 ;
        RECT 15.345 217.670 16.345 217.700 ;
        RECT 15.345 217.440 16.345 217.460 ;
        RECT 15.330 217.140 16.370 217.440 ;
        RECT 16.520 217.400 18.550 217.730 ;
        RECT 18.690 217.610 19.690 218.160 ;
        RECT 19.870 217.700 20.130 217.730 ;
        RECT 18.690 217.440 19.690 217.450 ;
        RECT 18.690 217.230 19.700 217.440 ;
        RECT 19.850 217.410 20.130 217.700 ;
        RECT 19.870 217.390 20.130 217.410 ;
        RECT 18.550 217.140 19.700 217.230 ;
        RECT 15.330 217.000 19.700 217.140 ;
        RECT 16.320 216.980 19.700 217.000 ;
        RECT 14.250 216.130 16.370 216.400 ;
        RECT 14.250 214.300 14.600 216.130 ;
        RECT 14.850 215.300 15.170 215.630 ;
        RECT 15.330 215.600 16.360 216.130 ;
        RECT 17.090 215.630 17.820 216.980 ;
        RECT 20.380 216.390 21.320 218.160 ;
        RECT 21.570 217.760 21.830 217.790 ;
        RECT 21.570 217.470 21.850 217.760 ;
        RECT 22.010 217.670 23.010 218.220 ;
        RECT 23.880 217.790 24.610 219.140 ;
        RECT 27.100 218.560 27.450 220.390 ;
        RECT 25.330 218.290 27.450 218.560 ;
        RECT 22.010 217.500 23.010 217.510 ;
        RECT 21.570 217.450 21.830 217.470 ;
        RECT 22.000 217.290 23.010 217.500 ;
        RECT 23.150 217.460 25.180 217.790 ;
        RECT 25.340 217.760 26.370 218.290 ;
        RECT 25.355 217.730 26.355 217.760 ;
        RECT 25.355 217.500 26.355 217.520 ;
        RECT 22.000 217.200 23.150 217.290 ;
        RECT 25.330 217.200 26.370 217.500 ;
        RECT 26.530 217.460 26.850 217.790 ;
        RECT 22.000 217.060 26.370 217.200 ;
        RECT 22.000 217.040 25.380 217.060 ;
        RECT 20.380 216.330 23.010 216.390 ;
        RECT 18.690 216.120 23.010 216.330 ;
        RECT 18.690 216.060 21.320 216.120 ;
        RECT 15.345 215.570 16.345 215.600 ;
        RECT 15.345 215.340 16.345 215.360 ;
        RECT 15.330 215.040 16.370 215.340 ;
        RECT 16.520 215.300 18.550 215.630 ;
        RECT 18.690 215.510 19.690 216.060 ;
        RECT 19.870 215.600 20.130 215.630 ;
        RECT 18.690 215.340 19.690 215.350 ;
        RECT 18.690 215.130 19.700 215.340 ;
        RECT 19.850 215.310 20.130 215.600 ;
        RECT 19.870 215.290 20.130 215.310 ;
        RECT 18.550 215.040 19.700 215.130 ;
        RECT 15.330 214.900 19.700 215.040 ;
        RECT 16.320 214.880 19.700 214.900 ;
        RECT 14.250 214.030 16.370 214.300 ;
        RECT 14.250 212.210 14.600 214.030 ;
        RECT 14.850 213.200 15.170 213.530 ;
        RECT 15.330 213.500 16.360 214.030 ;
        RECT 17.090 213.530 17.820 214.880 ;
        RECT 20.380 214.290 21.320 216.060 ;
        RECT 21.570 215.660 21.830 215.690 ;
        RECT 21.570 215.370 21.850 215.660 ;
        RECT 22.010 215.570 23.010 216.120 ;
        RECT 23.880 215.690 24.610 217.040 ;
        RECT 27.100 216.460 27.450 218.290 ;
        RECT 25.330 216.190 27.450 216.460 ;
        RECT 22.010 215.400 23.010 215.410 ;
        RECT 21.570 215.350 21.830 215.370 ;
        RECT 22.000 215.190 23.010 215.400 ;
        RECT 23.150 215.360 25.180 215.690 ;
        RECT 25.340 215.660 26.370 216.190 ;
        RECT 25.355 215.630 26.355 215.660 ;
        RECT 25.355 215.400 26.355 215.420 ;
        RECT 22.000 215.100 23.150 215.190 ;
        RECT 25.330 215.100 26.370 215.400 ;
        RECT 26.530 215.360 26.850 215.690 ;
        RECT 22.000 214.960 26.370 215.100 ;
        RECT 22.000 214.940 25.380 214.960 ;
        RECT 20.380 214.230 23.010 214.290 ;
        RECT 18.690 214.020 23.010 214.230 ;
        RECT 18.690 213.960 21.320 214.020 ;
        RECT 15.345 213.470 16.345 213.500 ;
        RECT 15.345 213.240 16.345 213.260 ;
        RECT 15.330 212.940 16.370 213.240 ;
        RECT 16.520 213.200 18.550 213.530 ;
        RECT 18.690 213.410 19.690 213.960 ;
        RECT 19.870 213.500 20.130 213.530 ;
        RECT 18.690 213.240 19.690 213.250 ;
        RECT 18.690 213.030 19.700 213.240 ;
        RECT 19.850 213.210 20.130 213.500 ;
        RECT 19.870 213.190 20.130 213.210 ;
        RECT 18.550 212.940 19.700 213.030 ;
        RECT 15.330 212.800 19.700 212.940 ;
        RECT 16.320 212.780 19.700 212.800 ;
        RECT 14.250 211.940 16.370 212.210 ;
        RECT 14.250 210.110 14.600 211.940 ;
        RECT 14.850 211.110 15.170 211.440 ;
        RECT 15.330 211.410 16.360 211.940 ;
        RECT 17.090 211.440 17.820 212.780 ;
        RECT 20.380 212.190 21.320 213.960 ;
        RECT 21.570 213.560 21.830 213.590 ;
        RECT 21.570 213.270 21.850 213.560 ;
        RECT 22.010 213.470 23.010 214.020 ;
        RECT 23.880 213.590 24.610 214.940 ;
        RECT 27.100 214.360 27.450 216.190 ;
        RECT 25.330 214.090 27.450 214.360 ;
        RECT 22.010 213.300 23.010 213.310 ;
        RECT 21.570 213.250 21.830 213.270 ;
        RECT 22.000 213.090 23.010 213.300 ;
        RECT 23.150 213.260 25.180 213.590 ;
        RECT 25.340 213.560 26.370 214.090 ;
        RECT 25.355 213.530 26.355 213.560 ;
        RECT 25.355 213.300 26.355 213.320 ;
        RECT 22.000 213.000 23.150 213.090 ;
        RECT 25.330 213.000 26.370 213.300 ;
        RECT 26.530 213.260 26.850 213.590 ;
        RECT 22.000 212.860 26.370 213.000 ;
        RECT 22.000 212.840 25.380 212.860 ;
        RECT 20.380 212.140 23.010 212.190 ;
        RECT 18.690 211.920 23.010 212.140 ;
        RECT 18.690 211.870 21.320 211.920 ;
        RECT 15.345 211.380 16.345 211.410 ;
        RECT 15.345 211.150 16.345 211.170 ;
        RECT 15.330 210.850 16.370 211.150 ;
        RECT 16.520 211.110 18.550 211.440 ;
        RECT 18.690 211.320 19.690 211.870 ;
        RECT 19.870 211.410 20.130 211.440 ;
        RECT 18.690 211.150 19.690 211.160 ;
        RECT 18.690 210.940 19.700 211.150 ;
        RECT 19.850 211.120 20.130 211.410 ;
        RECT 19.870 211.100 20.130 211.120 ;
        RECT 18.550 210.850 19.700 210.940 ;
        RECT 15.330 210.710 19.700 210.850 ;
        RECT 16.320 210.690 19.700 210.710 ;
        RECT 14.250 209.840 16.370 210.110 ;
        RECT 14.250 208.020 14.600 209.840 ;
        RECT 14.850 209.010 15.170 209.340 ;
        RECT 15.330 209.310 16.360 209.840 ;
        RECT 17.090 209.340 17.820 210.690 ;
        RECT 20.380 210.090 21.320 211.870 ;
        RECT 21.570 211.460 21.830 211.490 ;
        RECT 21.570 211.170 21.850 211.460 ;
        RECT 22.010 211.370 23.010 211.920 ;
        RECT 23.880 211.490 24.610 212.840 ;
        RECT 27.100 212.260 27.450 214.090 ;
        RECT 25.330 211.990 27.450 212.260 ;
        RECT 22.010 211.200 23.010 211.210 ;
        RECT 21.570 211.150 21.830 211.170 ;
        RECT 22.000 210.990 23.010 211.200 ;
        RECT 23.150 211.160 25.180 211.490 ;
        RECT 25.340 211.460 26.370 211.990 ;
        RECT 25.355 211.430 26.355 211.460 ;
        RECT 25.355 211.200 26.355 211.220 ;
        RECT 22.000 210.900 23.150 210.990 ;
        RECT 25.330 210.900 26.370 211.200 ;
        RECT 26.530 211.160 26.850 211.490 ;
        RECT 22.000 210.760 26.370 210.900 ;
        RECT 22.000 210.740 25.380 210.760 ;
        RECT 20.380 210.040 23.010 210.090 ;
        RECT 18.690 209.820 23.010 210.040 ;
        RECT 18.690 209.770 21.320 209.820 ;
        RECT 15.345 209.280 16.345 209.310 ;
        RECT 15.345 209.050 16.345 209.070 ;
        RECT 15.330 208.750 16.370 209.050 ;
        RECT 16.520 209.010 18.550 209.340 ;
        RECT 18.690 209.220 19.690 209.770 ;
        RECT 19.870 209.310 20.130 209.340 ;
        RECT 18.690 209.050 19.690 209.060 ;
        RECT 18.690 208.840 19.700 209.050 ;
        RECT 19.850 209.020 20.130 209.310 ;
        RECT 19.870 209.000 20.130 209.020 ;
        RECT 18.550 208.750 19.700 208.840 ;
        RECT 15.330 208.610 19.700 208.750 ;
        RECT 16.320 208.590 19.700 208.610 ;
        RECT 14.250 207.750 16.370 208.020 ;
        RECT 14.250 205.920 14.600 207.750 ;
        RECT 14.850 206.920 15.170 207.250 ;
        RECT 15.330 207.220 16.360 207.750 ;
        RECT 17.090 207.250 17.820 208.590 ;
        RECT 20.380 207.990 21.320 209.770 ;
        RECT 21.570 209.360 21.830 209.390 ;
        RECT 21.570 209.070 21.850 209.360 ;
        RECT 22.010 209.270 23.010 209.820 ;
        RECT 23.880 209.390 24.610 210.740 ;
        RECT 27.100 210.160 27.450 211.990 ;
        RECT 25.330 209.890 27.450 210.160 ;
        RECT 22.010 209.100 23.010 209.110 ;
        RECT 21.570 209.050 21.830 209.070 ;
        RECT 22.000 208.890 23.010 209.100 ;
        RECT 23.150 209.060 25.180 209.390 ;
        RECT 25.340 209.360 26.370 209.890 ;
        RECT 25.355 209.330 26.355 209.360 ;
        RECT 25.355 209.100 26.355 209.120 ;
        RECT 22.000 208.800 23.150 208.890 ;
        RECT 25.330 208.800 26.370 209.100 ;
        RECT 26.530 209.060 26.850 209.390 ;
        RECT 22.000 208.660 26.370 208.800 ;
        RECT 22.000 208.640 25.380 208.660 ;
        RECT 20.380 207.950 23.010 207.990 ;
        RECT 18.690 207.720 23.010 207.950 ;
        RECT 18.690 207.680 21.320 207.720 ;
        RECT 15.345 207.190 16.345 207.220 ;
        RECT 15.345 206.960 16.345 206.980 ;
        RECT 15.330 206.660 16.370 206.960 ;
        RECT 16.520 206.920 18.550 207.250 ;
        RECT 18.690 207.130 19.690 207.680 ;
        RECT 19.870 207.220 20.130 207.250 ;
        RECT 18.690 206.960 19.690 206.970 ;
        RECT 18.690 206.750 19.700 206.960 ;
        RECT 19.850 206.930 20.130 207.220 ;
        RECT 19.870 206.910 20.130 206.930 ;
        RECT 18.550 206.660 19.700 206.750 ;
        RECT 15.330 206.520 19.700 206.660 ;
        RECT 16.320 206.500 19.700 206.520 ;
        RECT 14.250 205.650 16.370 205.920 ;
        RECT 14.250 203.820 14.600 205.650 ;
        RECT 14.850 204.820 15.170 205.150 ;
        RECT 15.330 205.120 16.360 205.650 ;
        RECT 17.090 205.150 17.820 206.500 ;
        RECT 20.380 205.890 21.320 207.680 ;
        RECT 21.570 207.260 21.830 207.290 ;
        RECT 21.570 206.970 21.850 207.260 ;
        RECT 22.010 207.170 23.010 207.720 ;
        RECT 23.880 207.290 24.610 208.640 ;
        RECT 27.100 208.060 27.450 209.890 ;
        RECT 25.330 207.790 27.450 208.060 ;
        RECT 22.010 207.000 23.010 207.010 ;
        RECT 21.570 206.950 21.830 206.970 ;
        RECT 22.000 206.790 23.010 207.000 ;
        RECT 23.150 206.960 25.180 207.290 ;
        RECT 25.340 207.260 26.370 207.790 ;
        RECT 25.355 207.230 26.355 207.260 ;
        RECT 25.355 207.000 26.355 207.020 ;
        RECT 22.000 206.700 23.150 206.790 ;
        RECT 25.330 206.700 26.370 207.000 ;
        RECT 26.530 206.960 26.850 207.290 ;
        RECT 22.000 206.560 26.370 206.700 ;
        RECT 22.000 206.540 25.380 206.560 ;
        RECT 20.380 205.850 23.010 205.890 ;
        RECT 18.690 205.620 23.010 205.850 ;
        RECT 18.690 205.580 21.320 205.620 ;
        RECT 15.345 205.090 16.345 205.120 ;
        RECT 15.345 204.860 16.345 204.880 ;
        RECT 15.330 204.560 16.370 204.860 ;
        RECT 16.520 204.820 18.550 205.150 ;
        RECT 18.690 205.030 19.690 205.580 ;
        RECT 19.870 205.120 20.130 205.150 ;
        RECT 18.690 204.860 19.690 204.870 ;
        RECT 18.690 204.650 19.700 204.860 ;
        RECT 19.850 204.830 20.130 205.120 ;
        RECT 19.870 204.810 20.130 204.830 ;
        RECT 18.550 204.560 19.700 204.650 ;
        RECT 15.330 204.420 19.700 204.560 ;
        RECT 16.320 204.400 19.700 204.420 ;
        RECT 14.250 203.550 16.370 203.820 ;
        RECT 14.250 201.720 14.600 203.550 ;
        RECT 14.850 202.720 15.170 203.050 ;
        RECT 15.330 203.020 16.360 203.550 ;
        RECT 17.090 203.050 17.820 204.400 ;
        RECT 20.380 203.790 21.320 205.580 ;
        RECT 21.570 205.160 21.830 205.190 ;
        RECT 21.570 204.870 21.850 205.160 ;
        RECT 22.010 205.070 23.010 205.620 ;
        RECT 23.880 205.190 24.610 206.540 ;
        RECT 27.100 205.960 27.450 207.790 ;
        RECT 25.330 205.690 27.450 205.960 ;
        RECT 22.010 204.900 23.010 204.910 ;
        RECT 21.570 204.850 21.830 204.870 ;
        RECT 22.000 204.690 23.010 204.900 ;
        RECT 23.150 204.860 25.180 205.190 ;
        RECT 25.340 205.160 26.370 205.690 ;
        RECT 25.355 205.130 26.355 205.160 ;
        RECT 25.355 204.900 26.355 204.920 ;
        RECT 22.000 204.600 23.150 204.690 ;
        RECT 25.330 204.600 26.370 204.900 ;
        RECT 26.530 204.860 26.850 205.190 ;
        RECT 22.000 204.460 26.370 204.600 ;
        RECT 22.000 204.440 25.380 204.460 ;
        RECT 20.380 203.750 23.010 203.790 ;
        RECT 18.690 203.520 23.010 203.750 ;
        RECT 18.690 203.480 21.320 203.520 ;
        RECT 15.345 202.990 16.345 203.020 ;
        RECT 15.345 202.760 16.345 202.780 ;
        RECT 15.330 202.460 16.370 202.760 ;
        RECT 16.520 202.720 18.550 203.050 ;
        RECT 18.690 202.930 19.690 203.480 ;
        RECT 19.870 203.020 20.130 203.050 ;
        RECT 18.690 202.760 19.690 202.770 ;
        RECT 18.690 202.550 19.700 202.760 ;
        RECT 19.850 202.730 20.130 203.020 ;
        RECT 19.870 202.710 20.130 202.730 ;
        RECT 18.550 202.460 19.700 202.550 ;
        RECT 15.330 202.320 19.700 202.460 ;
        RECT 16.320 202.300 19.700 202.320 ;
        RECT 14.250 201.450 16.370 201.720 ;
        RECT 14.250 199.620 14.600 201.450 ;
        RECT 14.850 200.620 15.170 200.950 ;
        RECT 15.330 200.920 16.360 201.450 ;
        RECT 17.090 200.950 17.820 202.300 ;
        RECT 20.380 201.690 21.320 203.480 ;
        RECT 21.570 203.060 21.830 203.090 ;
        RECT 21.570 202.770 21.850 203.060 ;
        RECT 22.010 202.970 23.010 203.520 ;
        RECT 23.880 203.090 24.610 204.440 ;
        RECT 27.100 203.860 27.450 205.690 ;
        RECT 25.330 203.590 27.450 203.860 ;
        RECT 22.010 202.800 23.010 202.810 ;
        RECT 21.570 202.750 21.830 202.770 ;
        RECT 22.000 202.590 23.010 202.800 ;
        RECT 23.150 202.760 25.180 203.090 ;
        RECT 25.340 203.060 26.370 203.590 ;
        RECT 25.355 203.030 26.355 203.060 ;
        RECT 25.355 202.800 26.355 202.820 ;
        RECT 22.000 202.500 23.150 202.590 ;
        RECT 25.330 202.500 26.370 202.800 ;
        RECT 26.530 202.760 26.850 203.090 ;
        RECT 22.000 202.360 26.370 202.500 ;
        RECT 22.000 202.340 25.380 202.360 ;
        RECT 20.380 201.650 23.010 201.690 ;
        RECT 18.690 201.420 23.010 201.650 ;
        RECT 18.690 201.380 21.320 201.420 ;
        RECT 15.345 200.890 16.345 200.920 ;
        RECT 15.345 200.660 16.345 200.680 ;
        RECT 15.330 200.360 16.370 200.660 ;
        RECT 16.520 200.620 18.550 200.950 ;
        RECT 18.690 200.830 19.690 201.380 ;
        RECT 19.870 200.920 20.130 200.950 ;
        RECT 18.690 200.660 19.690 200.670 ;
        RECT 18.690 200.450 19.700 200.660 ;
        RECT 19.850 200.630 20.130 200.920 ;
        RECT 19.870 200.610 20.130 200.630 ;
        RECT 18.550 200.360 19.700 200.450 ;
        RECT 15.330 200.220 19.700 200.360 ;
        RECT 16.320 200.200 19.700 200.220 ;
        RECT 14.250 199.350 16.370 199.620 ;
        RECT 14.250 197.520 14.600 199.350 ;
        RECT 14.850 198.520 15.170 198.850 ;
        RECT 15.330 198.820 16.360 199.350 ;
        RECT 17.090 198.850 17.820 200.200 ;
        RECT 20.380 199.590 21.320 201.380 ;
        RECT 21.570 200.960 21.830 200.990 ;
        RECT 21.570 200.670 21.850 200.960 ;
        RECT 22.010 200.870 23.010 201.420 ;
        RECT 23.880 200.990 24.610 202.340 ;
        RECT 27.100 201.760 27.450 203.590 ;
        RECT 25.330 201.490 27.450 201.760 ;
        RECT 22.010 200.700 23.010 200.710 ;
        RECT 21.570 200.650 21.830 200.670 ;
        RECT 22.000 200.490 23.010 200.700 ;
        RECT 23.150 200.660 25.180 200.990 ;
        RECT 25.340 200.960 26.370 201.490 ;
        RECT 25.355 200.930 26.355 200.960 ;
        RECT 25.355 200.700 26.355 200.720 ;
        RECT 22.000 200.400 23.150 200.490 ;
        RECT 25.330 200.400 26.370 200.700 ;
        RECT 26.530 200.660 26.850 200.990 ;
        RECT 22.000 200.260 26.370 200.400 ;
        RECT 22.000 200.240 25.380 200.260 ;
        RECT 20.380 199.550 23.010 199.590 ;
        RECT 18.690 199.320 23.010 199.550 ;
        RECT 18.690 199.280 21.320 199.320 ;
        RECT 15.345 198.790 16.345 198.820 ;
        RECT 15.345 198.560 16.345 198.580 ;
        RECT 15.330 198.260 16.370 198.560 ;
        RECT 16.520 198.520 18.550 198.850 ;
        RECT 18.690 198.730 19.690 199.280 ;
        RECT 19.870 198.820 20.130 198.850 ;
        RECT 18.690 198.560 19.690 198.570 ;
        RECT 18.690 198.350 19.700 198.560 ;
        RECT 19.850 198.530 20.130 198.820 ;
        RECT 19.870 198.510 20.130 198.530 ;
        RECT 18.550 198.260 19.700 198.350 ;
        RECT 15.330 198.120 19.700 198.260 ;
        RECT 16.320 198.100 19.700 198.120 ;
        RECT 14.250 197.250 16.370 197.520 ;
        RECT 14.250 195.420 14.600 197.250 ;
        RECT 14.850 196.420 15.170 196.750 ;
        RECT 15.330 196.720 16.360 197.250 ;
        RECT 17.090 196.750 17.820 198.100 ;
        RECT 20.380 197.490 21.320 199.280 ;
        RECT 21.570 198.860 21.830 198.890 ;
        RECT 21.570 198.570 21.850 198.860 ;
        RECT 22.010 198.770 23.010 199.320 ;
        RECT 23.880 198.890 24.610 200.240 ;
        RECT 27.100 199.660 27.450 201.490 ;
        RECT 25.330 199.390 27.450 199.660 ;
        RECT 22.010 198.600 23.010 198.610 ;
        RECT 21.570 198.550 21.830 198.570 ;
        RECT 22.000 198.390 23.010 198.600 ;
        RECT 23.150 198.560 25.180 198.890 ;
        RECT 25.340 198.860 26.370 199.390 ;
        RECT 25.355 198.830 26.355 198.860 ;
        RECT 25.355 198.600 26.355 198.620 ;
        RECT 22.000 198.300 23.150 198.390 ;
        RECT 25.330 198.300 26.370 198.600 ;
        RECT 26.530 198.560 26.850 198.890 ;
        RECT 22.000 198.160 26.370 198.300 ;
        RECT 22.000 198.140 25.380 198.160 ;
        RECT 20.380 197.450 23.010 197.490 ;
        RECT 18.690 197.220 23.010 197.450 ;
        RECT 18.690 197.180 21.320 197.220 ;
        RECT 15.345 196.690 16.345 196.720 ;
        RECT 15.345 196.460 16.345 196.480 ;
        RECT 15.330 196.160 16.370 196.460 ;
        RECT 16.520 196.420 18.550 196.750 ;
        RECT 18.690 196.630 19.690 197.180 ;
        RECT 19.870 196.720 20.130 196.750 ;
        RECT 18.690 196.460 19.690 196.470 ;
        RECT 18.690 196.250 19.700 196.460 ;
        RECT 19.850 196.430 20.130 196.720 ;
        RECT 19.870 196.410 20.130 196.430 ;
        RECT 18.550 196.160 19.700 196.250 ;
        RECT 15.330 196.020 19.700 196.160 ;
        RECT 16.320 196.000 19.700 196.020 ;
        RECT 14.250 195.150 16.370 195.420 ;
        RECT 14.250 193.320 14.600 195.150 ;
        RECT 14.850 194.320 15.170 194.650 ;
        RECT 15.330 194.620 16.360 195.150 ;
        RECT 17.090 194.650 17.820 196.000 ;
        RECT 20.380 195.390 21.320 197.180 ;
        RECT 21.570 196.760 21.830 196.790 ;
        RECT 21.570 196.470 21.850 196.760 ;
        RECT 22.010 196.670 23.010 197.220 ;
        RECT 23.880 196.790 24.610 198.140 ;
        RECT 27.100 197.560 27.450 199.390 ;
        RECT 25.330 197.290 27.450 197.560 ;
        RECT 22.010 196.500 23.010 196.510 ;
        RECT 21.570 196.450 21.830 196.470 ;
        RECT 22.000 196.290 23.010 196.500 ;
        RECT 23.150 196.460 25.180 196.790 ;
        RECT 25.340 196.760 26.370 197.290 ;
        RECT 25.355 196.730 26.355 196.760 ;
        RECT 25.355 196.500 26.355 196.520 ;
        RECT 22.000 196.200 23.150 196.290 ;
        RECT 25.330 196.200 26.370 196.500 ;
        RECT 26.530 196.460 26.850 196.790 ;
        RECT 22.000 196.060 26.370 196.200 ;
        RECT 22.000 196.040 25.380 196.060 ;
        RECT 20.380 195.350 23.010 195.390 ;
        RECT 18.690 195.120 23.010 195.350 ;
        RECT 18.690 195.080 21.320 195.120 ;
        RECT 15.345 194.590 16.345 194.620 ;
        RECT 15.345 194.360 16.345 194.380 ;
        RECT 15.330 194.060 16.370 194.360 ;
        RECT 16.520 194.320 18.550 194.650 ;
        RECT 18.690 194.530 19.690 195.080 ;
        RECT 19.870 194.620 20.130 194.650 ;
        RECT 18.690 194.360 19.690 194.370 ;
        RECT 18.690 194.150 19.700 194.360 ;
        RECT 19.850 194.330 20.130 194.620 ;
        RECT 19.870 194.310 20.130 194.330 ;
        RECT 18.550 194.060 19.700 194.150 ;
        RECT 15.330 193.920 19.700 194.060 ;
        RECT 16.320 193.900 19.700 193.920 ;
        RECT 14.250 193.050 16.370 193.320 ;
        RECT 14.250 191.220 14.600 193.050 ;
        RECT 14.850 192.220 15.170 192.550 ;
        RECT 15.330 192.520 16.360 193.050 ;
        RECT 17.090 192.550 17.820 193.900 ;
        RECT 20.380 193.290 21.320 195.080 ;
        RECT 21.570 194.660 21.830 194.690 ;
        RECT 21.570 194.370 21.850 194.660 ;
        RECT 22.010 194.570 23.010 195.120 ;
        RECT 23.880 194.690 24.610 196.040 ;
        RECT 27.100 195.460 27.450 197.290 ;
        RECT 25.330 195.190 27.450 195.460 ;
        RECT 22.010 194.400 23.010 194.410 ;
        RECT 21.570 194.350 21.830 194.370 ;
        RECT 22.000 194.190 23.010 194.400 ;
        RECT 23.150 194.360 25.180 194.690 ;
        RECT 25.340 194.660 26.370 195.190 ;
        RECT 25.355 194.630 26.355 194.660 ;
        RECT 25.355 194.400 26.355 194.420 ;
        RECT 22.000 194.100 23.150 194.190 ;
        RECT 25.330 194.100 26.370 194.400 ;
        RECT 26.530 194.360 26.850 194.690 ;
        RECT 22.000 193.960 26.370 194.100 ;
        RECT 22.000 193.940 25.380 193.960 ;
        RECT 20.380 193.250 23.010 193.290 ;
        RECT 18.690 193.020 23.010 193.250 ;
        RECT 18.690 192.980 21.320 193.020 ;
        RECT 15.345 192.490 16.345 192.520 ;
        RECT 15.345 192.260 16.345 192.280 ;
        RECT 15.330 191.960 16.370 192.260 ;
        RECT 16.520 192.220 18.550 192.550 ;
        RECT 18.690 192.430 19.690 192.980 ;
        RECT 19.870 192.520 20.130 192.550 ;
        RECT 18.690 192.260 19.690 192.270 ;
        RECT 18.690 192.050 19.700 192.260 ;
        RECT 19.850 192.230 20.130 192.520 ;
        RECT 19.870 192.210 20.130 192.230 ;
        RECT 18.550 191.960 19.700 192.050 ;
        RECT 15.330 191.820 19.700 191.960 ;
        RECT 16.320 191.800 19.700 191.820 ;
        RECT 14.250 190.950 16.370 191.220 ;
        RECT 14.250 189.130 14.600 190.950 ;
        RECT 14.850 190.120 15.170 190.450 ;
        RECT 15.330 190.420 16.360 190.950 ;
        RECT 17.090 190.450 17.820 191.800 ;
        RECT 20.380 191.190 21.320 192.980 ;
        RECT 21.570 192.560 21.830 192.590 ;
        RECT 21.570 192.270 21.850 192.560 ;
        RECT 22.010 192.470 23.010 193.020 ;
        RECT 23.880 192.590 24.610 193.940 ;
        RECT 27.100 193.360 27.450 195.190 ;
        RECT 25.330 193.090 27.450 193.360 ;
        RECT 22.010 192.300 23.010 192.310 ;
        RECT 21.570 192.250 21.830 192.270 ;
        RECT 22.000 192.090 23.010 192.300 ;
        RECT 23.150 192.260 25.180 192.590 ;
        RECT 25.340 192.560 26.370 193.090 ;
        RECT 25.355 192.530 26.355 192.560 ;
        RECT 25.355 192.300 26.355 192.320 ;
        RECT 22.000 192.000 23.150 192.090 ;
        RECT 25.330 192.000 26.370 192.300 ;
        RECT 26.530 192.260 26.850 192.590 ;
        RECT 22.000 191.860 26.370 192.000 ;
        RECT 22.000 191.840 25.380 191.860 ;
        RECT 20.380 191.150 23.010 191.190 ;
        RECT 18.690 190.920 23.010 191.150 ;
        RECT 18.690 190.880 21.320 190.920 ;
        RECT 15.345 190.390 16.345 190.420 ;
        RECT 15.345 190.160 16.345 190.180 ;
        RECT 15.330 189.860 16.370 190.160 ;
        RECT 16.520 190.120 18.550 190.450 ;
        RECT 18.690 190.330 19.690 190.880 ;
        RECT 19.870 190.420 20.130 190.450 ;
        RECT 18.690 190.160 19.690 190.170 ;
        RECT 18.690 189.950 19.700 190.160 ;
        RECT 19.850 190.130 20.130 190.420 ;
        RECT 19.870 190.110 20.130 190.130 ;
        RECT 18.550 189.860 19.700 189.950 ;
        RECT 15.330 189.720 19.700 189.860 ;
        RECT 16.320 189.700 19.700 189.720 ;
        RECT 14.250 188.860 16.370 189.130 ;
        RECT 14.250 187.040 14.600 188.860 ;
        RECT 14.850 188.030 15.170 188.360 ;
        RECT 15.330 188.330 16.360 188.860 ;
        RECT 17.090 188.360 17.820 189.700 ;
        RECT 20.380 189.090 21.320 190.880 ;
        RECT 21.570 190.460 21.830 190.490 ;
        RECT 21.570 190.170 21.850 190.460 ;
        RECT 22.010 190.370 23.010 190.920 ;
        RECT 23.880 190.490 24.610 191.840 ;
        RECT 27.100 191.260 27.450 193.090 ;
        RECT 25.330 190.990 27.450 191.260 ;
        RECT 22.010 190.200 23.010 190.210 ;
        RECT 21.570 190.150 21.830 190.170 ;
        RECT 22.000 189.990 23.010 190.200 ;
        RECT 23.150 190.160 25.180 190.490 ;
        RECT 25.340 190.460 26.370 190.990 ;
        RECT 25.355 190.430 26.355 190.460 ;
        RECT 25.355 190.200 26.355 190.220 ;
        RECT 22.000 189.900 23.150 189.990 ;
        RECT 25.330 189.900 26.370 190.200 ;
        RECT 26.530 190.160 26.850 190.490 ;
        RECT 22.000 189.760 26.370 189.900 ;
        RECT 22.000 189.740 25.380 189.760 ;
        RECT 20.380 189.060 23.010 189.090 ;
        RECT 18.690 188.820 23.010 189.060 ;
        RECT 18.690 188.790 21.320 188.820 ;
        RECT 15.345 188.300 16.345 188.330 ;
        RECT 15.345 188.070 16.345 188.090 ;
        RECT 15.330 187.770 16.370 188.070 ;
        RECT 16.520 188.030 18.550 188.360 ;
        RECT 18.690 188.240 19.690 188.790 ;
        RECT 19.870 188.330 20.130 188.360 ;
        RECT 18.690 188.070 19.690 188.080 ;
        RECT 18.690 187.860 19.700 188.070 ;
        RECT 19.850 188.040 20.130 188.330 ;
        RECT 19.870 188.020 20.130 188.040 ;
        RECT 18.550 187.770 19.700 187.860 ;
        RECT 15.330 187.630 19.700 187.770 ;
        RECT 16.320 187.610 19.700 187.630 ;
        RECT 14.250 186.770 16.370 187.040 ;
        RECT 14.250 184.940 14.600 186.770 ;
        RECT 14.850 185.940 15.170 186.270 ;
        RECT 15.330 186.240 16.360 186.770 ;
        RECT 17.090 186.270 17.820 187.610 ;
        RECT 20.380 186.990 21.320 188.790 ;
        RECT 21.570 188.360 21.830 188.390 ;
        RECT 21.570 188.070 21.850 188.360 ;
        RECT 22.010 188.270 23.010 188.820 ;
        RECT 23.880 188.390 24.610 189.740 ;
        RECT 27.100 189.160 27.450 190.990 ;
        RECT 25.330 188.890 27.450 189.160 ;
        RECT 22.010 188.100 23.010 188.110 ;
        RECT 21.570 188.050 21.830 188.070 ;
        RECT 22.000 187.890 23.010 188.100 ;
        RECT 23.150 188.060 25.180 188.390 ;
        RECT 25.340 188.360 26.370 188.890 ;
        RECT 25.355 188.330 26.355 188.360 ;
        RECT 25.355 188.100 26.355 188.120 ;
        RECT 22.000 187.800 23.150 187.890 ;
        RECT 25.330 187.800 26.370 188.100 ;
        RECT 26.530 188.060 26.850 188.390 ;
        RECT 22.000 187.660 26.370 187.800 ;
        RECT 22.000 187.640 25.380 187.660 ;
        RECT 20.380 186.970 23.010 186.990 ;
        RECT 18.690 186.720 23.010 186.970 ;
        RECT 18.690 186.700 21.320 186.720 ;
        RECT 15.345 186.210 16.345 186.240 ;
        RECT 15.345 185.980 16.345 186.000 ;
        RECT 15.330 185.680 16.370 185.980 ;
        RECT 16.520 185.940 18.550 186.270 ;
        RECT 18.690 186.150 19.690 186.700 ;
        RECT 19.870 186.240 20.130 186.270 ;
        RECT 18.690 185.980 19.690 185.990 ;
        RECT 18.690 185.770 19.700 185.980 ;
        RECT 19.850 185.950 20.130 186.240 ;
        RECT 19.870 185.930 20.130 185.950 ;
        RECT 18.550 185.680 19.700 185.770 ;
        RECT 15.330 185.540 19.700 185.680 ;
        RECT 16.320 185.520 19.700 185.540 ;
        RECT 14.250 184.670 16.370 184.940 ;
        RECT 14.250 182.850 14.600 184.670 ;
        RECT 14.850 183.840 15.170 184.170 ;
        RECT 15.330 184.140 16.360 184.670 ;
        RECT 17.090 184.170 17.820 185.520 ;
        RECT 20.380 184.890 21.320 186.700 ;
        RECT 21.570 186.260 21.830 186.290 ;
        RECT 21.570 185.970 21.850 186.260 ;
        RECT 22.010 186.170 23.010 186.720 ;
        RECT 23.880 186.290 24.610 187.640 ;
        RECT 27.100 187.060 27.450 188.890 ;
        RECT 25.330 186.790 27.450 187.060 ;
        RECT 22.010 186.000 23.010 186.010 ;
        RECT 21.570 185.950 21.830 185.970 ;
        RECT 22.000 185.790 23.010 186.000 ;
        RECT 23.150 185.960 25.180 186.290 ;
        RECT 25.340 186.260 26.370 186.790 ;
        RECT 25.355 186.230 26.355 186.260 ;
        RECT 25.355 186.000 26.355 186.020 ;
        RECT 22.000 185.700 23.150 185.790 ;
        RECT 25.330 185.700 26.370 186.000 ;
        RECT 26.530 185.960 26.850 186.290 ;
        RECT 22.000 185.560 26.370 185.700 ;
        RECT 22.000 185.540 25.380 185.560 ;
        RECT 20.380 184.870 23.010 184.890 ;
        RECT 18.690 184.620 23.010 184.870 ;
        RECT 18.690 184.600 21.320 184.620 ;
        RECT 15.345 184.110 16.345 184.140 ;
        RECT 15.345 183.880 16.345 183.900 ;
        RECT 15.330 183.580 16.370 183.880 ;
        RECT 16.520 183.840 18.550 184.170 ;
        RECT 18.690 184.050 19.690 184.600 ;
        RECT 19.870 184.140 20.130 184.170 ;
        RECT 18.690 183.880 19.690 183.890 ;
        RECT 18.690 183.670 19.700 183.880 ;
        RECT 19.850 183.850 20.130 184.140 ;
        RECT 19.870 183.830 20.130 183.850 ;
        RECT 18.550 183.580 19.700 183.670 ;
        RECT 15.330 183.440 19.700 183.580 ;
        RECT 16.320 183.420 19.700 183.440 ;
        RECT 14.250 182.580 16.370 182.850 ;
        RECT 14.250 180.760 14.600 182.580 ;
        RECT 14.850 181.750 15.170 182.080 ;
        RECT 15.330 182.050 16.360 182.580 ;
        RECT 17.090 182.080 17.820 183.420 ;
        RECT 20.380 182.790 21.320 184.600 ;
        RECT 21.570 184.160 21.830 184.190 ;
        RECT 21.570 183.870 21.850 184.160 ;
        RECT 22.010 184.070 23.010 184.620 ;
        RECT 23.880 184.190 24.610 185.540 ;
        RECT 27.100 184.960 27.450 186.790 ;
        RECT 25.330 184.690 27.450 184.960 ;
        RECT 22.010 183.900 23.010 183.910 ;
        RECT 21.570 183.850 21.830 183.870 ;
        RECT 22.000 183.690 23.010 183.900 ;
        RECT 23.150 183.860 25.180 184.190 ;
        RECT 25.340 184.160 26.370 184.690 ;
        RECT 25.355 184.130 26.355 184.160 ;
        RECT 25.355 183.900 26.355 183.920 ;
        RECT 22.000 183.600 23.150 183.690 ;
        RECT 25.330 183.600 26.370 183.900 ;
        RECT 26.530 183.860 26.850 184.190 ;
        RECT 22.000 183.460 26.370 183.600 ;
        RECT 22.000 183.440 25.380 183.460 ;
        RECT 20.380 182.780 23.010 182.790 ;
        RECT 18.690 182.520 23.010 182.780 ;
        RECT 18.690 182.510 21.320 182.520 ;
        RECT 15.345 182.020 16.345 182.050 ;
        RECT 15.345 181.790 16.345 181.810 ;
        RECT 15.330 181.490 16.370 181.790 ;
        RECT 16.520 181.750 18.550 182.080 ;
        RECT 18.690 181.960 19.690 182.510 ;
        RECT 19.870 182.050 20.130 182.080 ;
        RECT 18.690 181.790 19.690 181.800 ;
        RECT 18.690 181.580 19.700 181.790 ;
        RECT 19.850 181.760 20.130 182.050 ;
        RECT 19.870 181.740 20.130 181.760 ;
        RECT 18.550 181.490 19.700 181.580 ;
        RECT 15.330 181.350 19.700 181.490 ;
        RECT 16.320 181.330 19.700 181.350 ;
        RECT 14.250 180.490 16.370 180.760 ;
        RECT 14.250 178.660 14.600 180.490 ;
        RECT 14.850 179.660 15.170 179.990 ;
        RECT 15.330 179.960 16.360 180.490 ;
        RECT 17.090 179.990 17.820 181.330 ;
        RECT 20.380 180.690 21.320 182.510 ;
        RECT 21.570 182.060 21.830 182.090 ;
        RECT 21.570 181.770 21.850 182.060 ;
        RECT 22.010 181.970 23.010 182.520 ;
        RECT 23.880 182.090 24.610 183.440 ;
        RECT 27.100 182.860 27.450 184.690 ;
        RECT 25.330 182.590 27.450 182.860 ;
        RECT 22.010 181.800 23.010 181.810 ;
        RECT 21.570 181.750 21.830 181.770 ;
        RECT 22.000 181.590 23.010 181.800 ;
        RECT 23.150 181.760 25.180 182.090 ;
        RECT 25.340 182.060 26.370 182.590 ;
        RECT 25.355 182.030 26.355 182.060 ;
        RECT 25.355 181.800 26.355 181.820 ;
        RECT 22.000 181.500 23.150 181.590 ;
        RECT 25.330 181.500 26.370 181.800 ;
        RECT 26.530 181.760 26.850 182.090 ;
        RECT 22.000 181.360 26.370 181.500 ;
        RECT 22.000 181.340 25.380 181.360 ;
        RECT 18.690 180.420 23.010 180.690 ;
        RECT 15.345 179.930 16.345 179.960 ;
        RECT 15.345 179.700 16.345 179.720 ;
        RECT 15.330 179.400 16.370 179.700 ;
        RECT 16.520 179.660 18.550 179.990 ;
        RECT 18.690 179.870 19.690 180.420 ;
        RECT 19.870 179.960 20.130 179.990 ;
        RECT 18.690 179.700 19.690 179.710 ;
        RECT 18.690 179.490 19.700 179.700 ;
        RECT 19.850 179.670 20.130 179.960 ;
        RECT 19.870 179.650 20.130 179.670 ;
        RECT 18.550 179.400 19.700 179.490 ;
        RECT 15.330 179.260 19.700 179.400 ;
        RECT 16.320 179.240 19.700 179.260 ;
        RECT 14.250 178.390 16.370 178.660 ;
        RECT 14.250 176.560 14.600 178.390 ;
        RECT 14.850 177.560 15.170 177.890 ;
        RECT 15.330 177.860 16.360 178.390 ;
        RECT 17.090 177.890 17.820 179.240 ;
        RECT 20.380 178.590 21.320 180.420 ;
        RECT 21.570 179.960 21.830 179.990 ;
        RECT 21.570 179.670 21.850 179.960 ;
        RECT 22.010 179.870 23.010 180.420 ;
        RECT 23.880 179.990 24.610 181.340 ;
        RECT 27.100 180.760 27.450 182.590 ;
        RECT 25.330 180.490 27.450 180.760 ;
        RECT 22.010 179.700 23.010 179.710 ;
        RECT 21.570 179.650 21.830 179.670 ;
        RECT 22.000 179.490 23.010 179.700 ;
        RECT 23.150 179.660 25.180 179.990 ;
        RECT 25.340 179.960 26.370 180.490 ;
        RECT 25.355 179.930 26.355 179.960 ;
        RECT 25.355 179.700 26.355 179.720 ;
        RECT 22.000 179.400 23.150 179.490 ;
        RECT 25.330 179.400 26.370 179.700 ;
        RECT 26.530 179.660 26.850 179.990 ;
        RECT 22.000 179.260 26.370 179.400 ;
        RECT 22.000 179.240 25.380 179.260 ;
        RECT 18.690 178.320 23.010 178.590 ;
        RECT 15.345 177.830 16.345 177.860 ;
        RECT 15.345 177.600 16.345 177.620 ;
        RECT 15.330 177.300 16.370 177.600 ;
        RECT 16.520 177.560 18.550 177.890 ;
        RECT 18.690 177.770 19.690 178.320 ;
        RECT 19.870 177.860 20.130 177.890 ;
        RECT 18.690 177.600 19.690 177.610 ;
        RECT 18.690 177.390 19.700 177.600 ;
        RECT 19.850 177.570 20.130 177.860 ;
        RECT 19.870 177.550 20.130 177.570 ;
        RECT 18.550 177.300 19.700 177.390 ;
        RECT 15.330 177.160 19.700 177.300 ;
        RECT 16.320 177.140 19.700 177.160 ;
        RECT 14.250 176.290 16.370 176.560 ;
        RECT 14.250 174.460 14.600 176.290 ;
        RECT 14.850 175.460 15.170 175.790 ;
        RECT 15.330 175.760 16.360 176.290 ;
        RECT 17.090 175.790 17.820 177.140 ;
        RECT 20.380 176.490 21.320 178.320 ;
        RECT 21.570 177.860 21.830 177.890 ;
        RECT 21.570 177.570 21.850 177.860 ;
        RECT 22.010 177.770 23.010 178.320 ;
        RECT 23.880 177.890 24.610 179.240 ;
        RECT 27.100 178.660 27.450 180.490 ;
        RECT 25.330 178.390 27.450 178.660 ;
        RECT 22.010 177.600 23.010 177.610 ;
        RECT 21.570 177.550 21.830 177.570 ;
        RECT 22.000 177.390 23.010 177.600 ;
        RECT 23.150 177.560 25.180 177.890 ;
        RECT 25.340 177.860 26.370 178.390 ;
        RECT 25.355 177.830 26.355 177.860 ;
        RECT 25.355 177.600 26.355 177.620 ;
        RECT 22.000 177.300 23.150 177.390 ;
        RECT 25.330 177.300 26.370 177.600 ;
        RECT 26.530 177.560 26.850 177.890 ;
        RECT 22.000 177.160 26.370 177.300 ;
        RECT 22.000 177.140 25.380 177.160 ;
        RECT 18.690 176.220 23.010 176.490 ;
        RECT 15.345 175.730 16.345 175.760 ;
        RECT 15.345 175.500 16.345 175.520 ;
        RECT 15.330 175.200 16.370 175.500 ;
        RECT 16.520 175.460 18.550 175.790 ;
        RECT 18.690 175.670 19.690 176.220 ;
        RECT 19.870 175.760 20.130 175.790 ;
        RECT 18.690 175.500 19.690 175.510 ;
        RECT 18.690 175.290 19.700 175.500 ;
        RECT 19.850 175.470 20.130 175.760 ;
        RECT 19.870 175.450 20.130 175.470 ;
        RECT 18.550 175.200 19.700 175.290 ;
        RECT 15.330 175.060 19.700 175.200 ;
        RECT 16.320 175.040 19.700 175.060 ;
        RECT 14.250 174.190 16.370 174.460 ;
        RECT 14.250 172.360 14.600 174.190 ;
        RECT 14.850 173.360 15.170 173.690 ;
        RECT 15.330 173.660 16.360 174.190 ;
        RECT 17.090 173.690 17.820 175.040 ;
        RECT 20.380 174.390 21.320 176.220 ;
        RECT 21.570 175.760 21.830 175.790 ;
        RECT 21.570 175.470 21.850 175.760 ;
        RECT 22.010 175.670 23.010 176.220 ;
        RECT 23.880 175.790 24.610 177.140 ;
        RECT 27.100 176.560 27.450 178.390 ;
        RECT 25.330 176.290 27.450 176.560 ;
        RECT 22.010 175.500 23.010 175.510 ;
        RECT 21.570 175.450 21.830 175.470 ;
        RECT 22.000 175.290 23.010 175.500 ;
        RECT 23.150 175.460 25.180 175.790 ;
        RECT 25.340 175.760 26.370 176.290 ;
        RECT 25.355 175.730 26.355 175.760 ;
        RECT 25.355 175.500 26.355 175.520 ;
        RECT 22.000 175.200 23.150 175.290 ;
        RECT 25.330 175.200 26.370 175.500 ;
        RECT 26.530 175.460 26.850 175.790 ;
        RECT 22.000 175.060 26.370 175.200 ;
        RECT 22.000 175.040 25.380 175.060 ;
        RECT 18.690 174.120 23.010 174.390 ;
        RECT 15.345 173.630 16.345 173.660 ;
        RECT 15.345 173.400 16.345 173.420 ;
        RECT 15.330 173.100 16.370 173.400 ;
        RECT 16.520 173.360 18.550 173.690 ;
        RECT 18.690 173.570 19.690 174.120 ;
        RECT 19.870 173.660 20.130 173.690 ;
        RECT 18.690 173.400 19.690 173.410 ;
        RECT 18.690 173.190 19.700 173.400 ;
        RECT 19.850 173.370 20.130 173.660 ;
        RECT 19.870 173.350 20.130 173.370 ;
        RECT 18.550 173.100 19.700 173.190 ;
        RECT 15.330 172.960 19.700 173.100 ;
        RECT 16.320 172.940 19.700 172.960 ;
        RECT 14.250 172.090 16.370 172.360 ;
        RECT 14.250 170.260 14.600 172.090 ;
        RECT 14.850 171.260 15.170 171.590 ;
        RECT 15.330 171.560 16.360 172.090 ;
        RECT 17.090 171.590 17.820 172.940 ;
        RECT 20.380 172.290 21.320 174.120 ;
        RECT 21.570 173.660 21.830 173.690 ;
        RECT 21.570 173.370 21.850 173.660 ;
        RECT 22.010 173.570 23.010 174.120 ;
        RECT 23.880 173.690 24.610 175.040 ;
        RECT 27.100 174.460 27.450 176.290 ;
        RECT 25.330 174.190 27.450 174.460 ;
        RECT 22.010 173.400 23.010 173.410 ;
        RECT 21.570 173.350 21.830 173.370 ;
        RECT 22.000 173.190 23.010 173.400 ;
        RECT 23.150 173.360 25.180 173.690 ;
        RECT 25.340 173.660 26.370 174.190 ;
        RECT 25.355 173.630 26.355 173.660 ;
        RECT 25.355 173.400 26.355 173.420 ;
        RECT 22.000 173.100 23.150 173.190 ;
        RECT 25.330 173.100 26.370 173.400 ;
        RECT 26.530 173.360 26.850 173.690 ;
        RECT 22.000 172.960 26.370 173.100 ;
        RECT 22.000 172.940 25.380 172.960 ;
        RECT 18.690 172.020 23.010 172.290 ;
        RECT 15.345 171.530 16.345 171.560 ;
        RECT 15.345 171.300 16.345 171.320 ;
        RECT 15.330 171.000 16.370 171.300 ;
        RECT 16.520 171.260 18.550 171.590 ;
        RECT 18.690 171.470 19.690 172.020 ;
        RECT 19.870 171.560 20.130 171.590 ;
        RECT 18.690 171.300 19.690 171.310 ;
        RECT 18.690 171.090 19.700 171.300 ;
        RECT 19.850 171.270 20.130 171.560 ;
        RECT 19.870 171.250 20.130 171.270 ;
        RECT 18.550 171.000 19.700 171.090 ;
        RECT 15.330 170.860 19.700 171.000 ;
        RECT 16.320 170.840 19.700 170.860 ;
        RECT 14.250 169.990 16.370 170.260 ;
        RECT 14.250 168.160 14.600 169.990 ;
        RECT 14.850 169.160 15.170 169.490 ;
        RECT 15.330 169.460 16.360 169.990 ;
        RECT 17.090 169.490 17.820 170.840 ;
        RECT 20.380 170.190 21.320 172.020 ;
        RECT 21.570 171.560 21.830 171.590 ;
        RECT 21.570 171.270 21.850 171.560 ;
        RECT 22.010 171.470 23.010 172.020 ;
        RECT 23.880 171.590 24.610 172.940 ;
        RECT 27.100 172.360 27.450 174.190 ;
        RECT 25.330 172.090 27.450 172.360 ;
        RECT 22.010 171.300 23.010 171.310 ;
        RECT 21.570 171.250 21.830 171.270 ;
        RECT 22.000 171.090 23.010 171.300 ;
        RECT 23.150 171.260 25.180 171.590 ;
        RECT 25.340 171.560 26.370 172.090 ;
        RECT 25.355 171.530 26.355 171.560 ;
        RECT 25.355 171.300 26.355 171.320 ;
        RECT 22.000 171.000 23.150 171.090 ;
        RECT 25.330 171.000 26.370 171.300 ;
        RECT 26.530 171.260 26.850 171.590 ;
        RECT 22.000 170.860 26.370 171.000 ;
        RECT 22.000 170.840 25.380 170.860 ;
        RECT 18.690 169.920 23.010 170.190 ;
        RECT 15.345 169.430 16.345 169.460 ;
        RECT 15.345 169.200 16.345 169.220 ;
        RECT 15.330 168.900 16.370 169.200 ;
        RECT 16.520 169.160 18.550 169.490 ;
        RECT 18.690 169.370 19.690 169.920 ;
        RECT 19.870 169.460 20.130 169.490 ;
        RECT 18.690 169.200 19.690 169.210 ;
        RECT 18.690 168.990 19.700 169.200 ;
        RECT 19.850 169.170 20.130 169.460 ;
        RECT 19.870 169.150 20.130 169.170 ;
        RECT 18.550 168.900 19.700 168.990 ;
        RECT 15.330 168.760 19.700 168.900 ;
        RECT 16.320 168.740 19.700 168.760 ;
        RECT 14.250 167.890 16.370 168.160 ;
        RECT 14.250 166.060 14.600 167.890 ;
        RECT 14.850 167.060 15.170 167.390 ;
        RECT 15.330 167.360 16.360 167.890 ;
        RECT 17.090 167.390 17.820 168.740 ;
        RECT 20.380 168.090 21.320 169.920 ;
        RECT 21.570 169.460 21.830 169.490 ;
        RECT 21.570 169.170 21.850 169.460 ;
        RECT 22.010 169.370 23.010 169.920 ;
        RECT 23.880 169.490 24.610 170.840 ;
        RECT 27.100 170.260 27.450 172.090 ;
        RECT 25.330 169.990 27.450 170.260 ;
        RECT 22.010 169.200 23.010 169.210 ;
        RECT 21.570 169.150 21.830 169.170 ;
        RECT 22.000 168.990 23.010 169.200 ;
        RECT 23.150 169.160 25.180 169.490 ;
        RECT 25.340 169.460 26.370 169.990 ;
        RECT 25.355 169.430 26.355 169.460 ;
        RECT 25.355 169.200 26.355 169.220 ;
        RECT 22.000 168.900 23.150 168.990 ;
        RECT 25.330 168.900 26.370 169.200 ;
        RECT 26.530 169.160 26.850 169.490 ;
        RECT 22.000 168.760 26.370 168.900 ;
        RECT 22.000 168.740 25.380 168.760 ;
        RECT 18.690 167.820 23.010 168.090 ;
        RECT 15.345 167.330 16.345 167.360 ;
        RECT 15.345 167.100 16.345 167.120 ;
        RECT 15.330 166.800 16.370 167.100 ;
        RECT 16.520 167.060 18.550 167.390 ;
        RECT 18.690 167.270 19.690 167.820 ;
        RECT 19.870 167.360 20.130 167.390 ;
        RECT 18.690 167.100 19.690 167.110 ;
        RECT 18.690 166.890 19.700 167.100 ;
        RECT 19.850 167.070 20.130 167.360 ;
        RECT 19.870 167.050 20.130 167.070 ;
        RECT 18.550 166.800 19.700 166.890 ;
        RECT 15.330 166.660 19.700 166.800 ;
        RECT 16.320 166.640 19.700 166.660 ;
        RECT 14.250 165.790 16.370 166.060 ;
        RECT 14.250 163.960 14.600 165.790 ;
        RECT 14.850 164.960 15.170 165.290 ;
        RECT 15.330 165.260 16.360 165.790 ;
        RECT 17.090 165.290 17.820 166.640 ;
        RECT 20.380 165.990 21.320 167.820 ;
        RECT 21.570 167.360 21.830 167.390 ;
        RECT 21.570 167.070 21.850 167.360 ;
        RECT 22.010 167.270 23.010 167.820 ;
        RECT 23.880 167.390 24.610 168.740 ;
        RECT 27.100 168.160 27.450 169.990 ;
        RECT 25.330 167.890 27.450 168.160 ;
        RECT 22.010 167.100 23.010 167.110 ;
        RECT 21.570 167.050 21.830 167.070 ;
        RECT 22.000 166.890 23.010 167.100 ;
        RECT 23.150 167.060 25.180 167.390 ;
        RECT 25.340 167.360 26.370 167.890 ;
        RECT 25.355 167.330 26.355 167.360 ;
        RECT 25.355 167.100 26.355 167.120 ;
        RECT 22.000 166.800 23.150 166.890 ;
        RECT 25.330 166.800 26.370 167.100 ;
        RECT 26.530 167.060 26.850 167.390 ;
        RECT 22.000 166.660 26.370 166.800 ;
        RECT 22.000 166.640 25.380 166.660 ;
        RECT 18.690 165.720 23.010 165.990 ;
        RECT 15.345 165.230 16.345 165.260 ;
        RECT 15.345 165.000 16.345 165.020 ;
        RECT 15.330 164.700 16.370 165.000 ;
        RECT 16.520 164.960 18.550 165.290 ;
        RECT 18.690 165.170 19.690 165.720 ;
        RECT 19.870 165.260 20.130 165.290 ;
        RECT 18.690 165.000 19.690 165.010 ;
        RECT 18.690 164.790 19.700 165.000 ;
        RECT 19.850 164.970 20.130 165.260 ;
        RECT 19.870 164.950 20.130 164.970 ;
        RECT 18.550 164.700 19.700 164.790 ;
        RECT 15.330 164.560 19.700 164.700 ;
        RECT 16.320 164.540 19.700 164.560 ;
        RECT 14.250 163.690 16.370 163.960 ;
        RECT 14.250 161.860 14.600 163.690 ;
        RECT 14.850 162.860 15.170 163.190 ;
        RECT 15.330 163.160 16.360 163.690 ;
        RECT 17.090 163.190 17.820 164.540 ;
        RECT 20.380 163.890 21.320 165.720 ;
        RECT 21.570 165.260 21.830 165.290 ;
        RECT 21.570 164.970 21.850 165.260 ;
        RECT 22.010 165.170 23.010 165.720 ;
        RECT 23.880 165.290 24.610 166.640 ;
        RECT 27.100 166.060 27.450 167.890 ;
        RECT 25.330 165.790 27.450 166.060 ;
        RECT 22.010 165.000 23.010 165.010 ;
        RECT 21.570 164.950 21.830 164.970 ;
        RECT 22.000 164.790 23.010 165.000 ;
        RECT 23.150 164.960 25.180 165.290 ;
        RECT 25.340 165.260 26.370 165.790 ;
        RECT 25.355 165.230 26.355 165.260 ;
        RECT 25.355 165.000 26.355 165.020 ;
        RECT 22.000 164.700 23.150 164.790 ;
        RECT 25.330 164.700 26.370 165.000 ;
        RECT 26.530 164.960 26.850 165.290 ;
        RECT 22.000 164.560 26.370 164.700 ;
        RECT 22.000 164.540 25.380 164.560 ;
        RECT 18.690 163.620 23.010 163.890 ;
        RECT 15.345 163.130 16.345 163.160 ;
        RECT 15.345 162.900 16.345 162.920 ;
        RECT 15.330 162.600 16.370 162.900 ;
        RECT 16.520 162.860 18.550 163.190 ;
        RECT 18.690 163.070 19.690 163.620 ;
        RECT 19.870 163.160 20.130 163.190 ;
        RECT 18.690 162.900 19.690 162.910 ;
        RECT 18.690 162.690 19.700 162.900 ;
        RECT 19.850 162.870 20.130 163.160 ;
        RECT 19.870 162.850 20.130 162.870 ;
        RECT 18.550 162.600 19.700 162.690 ;
        RECT 15.330 162.460 19.700 162.600 ;
        RECT 16.320 162.440 19.700 162.460 ;
        RECT 14.250 161.590 16.370 161.860 ;
        RECT 14.250 159.760 14.600 161.590 ;
        RECT 14.850 160.760 15.170 161.090 ;
        RECT 15.330 161.060 16.360 161.590 ;
        RECT 17.090 161.090 17.820 162.440 ;
        RECT 20.380 161.790 21.320 163.620 ;
        RECT 21.570 163.160 21.830 163.190 ;
        RECT 21.570 162.870 21.850 163.160 ;
        RECT 22.010 163.070 23.010 163.620 ;
        RECT 23.880 163.190 24.610 164.540 ;
        RECT 27.100 163.960 27.450 165.790 ;
        RECT 25.330 163.690 27.450 163.960 ;
        RECT 22.010 162.900 23.010 162.910 ;
        RECT 21.570 162.850 21.830 162.870 ;
        RECT 22.000 162.690 23.010 162.900 ;
        RECT 23.150 162.860 25.180 163.190 ;
        RECT 25.340 163.160 26.370 163.690 ;
        RECT 25.355 163.130 26.355 163.160 ;
        RECT 25.355 162.900 26.355 162.920 ;
        RECT 22.000 162.600 23.150 162.690 ;
        RECT 25.330 162.600 26.370 162.900 ;
        RECT 26.530 162.860 26.850 163.190 ;
        RECT 22.000 162.460 26.370 162.600 ;
        RECT 22.000 162.440 25.380 162.460 ;
        RECT 18.690 161.520 23.010 161.790 ;
        RECT 15.345 161.030 16.345 161.060 ;
        RECT 15.345 160.800 16.345 160.820 ;
        RECT 15.330 160.500 16.370 160.800 ;
        RECT 16.520 160.760 18.550 161.090 ;
        RECT 18.690 160.970 19.690 161.520 ;
        RECT 19.870 161.060 20.130 161.090 ;
        RECT 18.690 160.800 19.690 160.810 ;
        RECT 18.690 160.590 19.700 160.800 ;
        RECT 19.850 160.770 20.130 161.060 ;
        RECT 19.870 160.750 20.130 160.770 ;
        RECT 18.550 160.500 19.700 160.590 ;
        RECT 15.330 160.360 19.700 160.500 ;
        RECT 16.320 160.340 19.700 160.360 ;
        RECT 14.250 159.490 16.370 159.760 ;
        RECT 14.250 157.660 14.600 159.490 ;
        RECT 14.850 158.660 15.170 158.990 ;
        RECT 15.330 158.960 16.360 159.490 ;
        RECT 17.090 158.990 17.820 160.340 ;
        RECT 20.380 159.690 21.320 161.520 ;
        RECT 21.570 161.060 21.830 161.090 ;
        RECT 21.570 160.770 21.850 161.060 ;
        RECT 22.010 160.970 23.010 161.520 ;
        RECT 23.880 161.090 24.610 162.440 ;
        RECT 27.100 161.860 27.450 163.690 ;
        RECT 25.330 161.590 27.450 161.860 ;
        RECT 22.010 160.800 23.010 160.810 ;
        RECT 21.570 160.750 21.830 160.770 ;
        RECT 22.000 160.590 23.010 160.800 ;
        RECT 23.150 160.760 25.180 161.090 ;
        RECT 25.340 161.060 26.370 161.590 ;
        RECT 25.355 161.030 26.355 161.060 ;
        RECT 25.355 160.800 26.355 160.820 ;
        RECT 22.000 160.500 23.150 160.590 ;
        RECT 25.330 160.500 26.370 160.800 ;
        RECT 26.530 160.760 26.850 161.090 ;
        RECT 22.000 160.360 26.370 160.500 ;
        RECT 22.000 160.340 25.380 160.360 ;
        RECT 18.690 159.420 23.010 159.690 ;
        RECT 15.345 158.930 16.345 158.960 ;
        RECT 15.345 158.700 16.345 158.720 ;
        RECT 15.330 158.400 16.370 158.700 ;
        RECT 16.520 158.660 18.550 158.990 ;
        RECT 18.690 158.870 19.690 159.420 ;
        RECT 19.870 158.960 20.130 158.990 ;
        RECT 18.690 158.700 19.690 158.710 ;
        RECT 18.690 158.490 19.700 158.700 ;
        RECT 19.850 158.670 20.130 158.960 ;
        RECT 19.870 158.650 20.130 158.670 ;
        RECT 18.550 158.400 19.700 158.490 ;
        RECT 15.330 158.260 19.700 158.400 ;
        RECT 16.320 158.240 19.700 158.260 ;
        RECT 14.250 157.390 16.370 157.660 ;
        RECT 14.250 155.560 14.600 157.390 ;
        RECT 14.850 156.560 15.170 156.890 ;
        RECT 15.330 156.860 16.360 157.390 ;
        RECT 17.090 156.890 17.820 158.240 ;
        RECT 20.380 157.590 21.320 159.420 ;
        RECT 21.570 158.960 21.830 158.990 ;
        RECT 21.570 158.670 21.850 158.960 ;
        RECT 22.010 158.870 23.010 159.420 ;
        RECT 23.880 158.990 24.610 160.340 ;
        RECT 27.100 159.760 27.450 161.590 ;
        RECT 25.330 159.490 27.450 159.760 ;
        RECT 22.010 158.700 23.010 158.710 ;
        RECT 21.570 158.650 21.830 158.670 ;
        RECT 22.000 158.490 23.010 158.700 ;
        RECT 23.150 158.660 25.180 158.990 ;
        RECT 25.340 158.960 26.370 159.490 ;
        RECT 25.355 158.930 26.355 158.960 ;
        RECT 25.355 158.700 26.355 158.720 ;
        RECT 22.000 158.400 23.150 158.490 ;
        RECT 25.330 158.400 26.370 158.700 ;
        RECT 26.530 158.660 26.850 158.990 ;
        RECT 22.000 158.260 26.370 158.400 ;
        RECT 22.000 158.240 25.380 158.260 ;
        RECT 18.690 157.320 23.010 157.590 ;
        RECT 15.345 156.830 16.345 156.860 ;
        RECT 15.345 156.600 16.345 156.620 ;
        RECT 15.330 156.300 16.370 156.600 ;
        RECT 16.520 156.560 18.550 156.890 ;
        RECT 18.690 156.770 19.690 157.320 ;
        RECT 19.870 156.860 20.130 156.890 ;
        RECT 18.690 156.600 19.690 156.610 ;
        RECT 18.690 156.390 19.700 156.600 ;
        RECT 19.850 156.570 20.130 156.860 ;
        RECT 19.870 156.550 20.130 156.570 ;
        RECT 18.550 156.300 19.700 156.390 ;
        RECT 15.330 156.160 19.700 156.300 ;
        RECT 16.320 156.140 19.700 156.160 ;
        RECT 14.250 155.290 16.370 155.560 ;
        RECT 14.250 153.460 14.600 155.290 ;
        RECT 14.850 154.460 15.170 154.790 ;
        RECT 15.330 154.760 16.360 155.290 ;
        RECT 17.090 154.790 17.820 156.140 ;
        RECT 20.380 155.490 21.320 157.320 ;
        RECT 21.570 156.860 21.830 156.890 ;
        RECT 21.570 156.570 21.850 156.860 ;
        RECT 22.010 156.770 23.010 157.320 ;
        RECT 23.880 156.890 24.610 158.240 ;
        RECT 27.100 157.660 27.450 159.490 ;
        RECT 25.330 157.390 27.450 157.660 ;
        RECT 22.010 156.600 23.010 156.610 ;
        RECT 21.570 156.550 21.830 156.570 ;
        RECT 22.000 156.390 23.010 156.600 ;
        RECT 23.150 156.560 25.180 156.890 ;
        RECT 25.340 156.860 26.370 157.390 ;
        RECT 25.355 156.830 26.355 156.860 ;
        RECT 25.355 156.600 26.355 156.620 ;
        RECT 22.000 156.300 23.150 156.390 ;
        RECT 25.330 156.300 26.370 156.600 ;
        RECT 26.530 156.560 26.850 156.890 ;
        RECT 22.000 156.160 26.370 156.300 ;
        RECT 22.000 156.140 25.380 156.160 ;
        RECT 18.690 155.220 23.010 155.490 ;
        RECT 15.345 154.730 16.345 154.760 ;
        RECT 15.345 154.500 16.345 154.520 ;
        RECT 15.330 154.200 16.370 154.500 ;
        RECT 16.520 154.460 18.550 154.790 ;
        RECT 18.690 154.670 19.690 155.220 ;
        RECT 19.870 154.760 20.130 154.790 ;
        RECT 18.690 154.500 19.690 154.510 ;
        RECT 18.690 154.290 19.700 154.500 ;
        RECT 19.850 154.470 20.130 154.760 ;
        RECT 19.870 154.450 20.130 154.470 ;
        RECT 18.550 154.200 19.700 154.290 ;
        RECT 15.330 154.060 19.700 154.200 ;
        RECT 16.320 154.040 19.700 154.060 ;
        RECT 14.250 153.190 16.370 153.460 ;
        RECT 14.250 151.360 14.600 153.190 ;
        RECT 14.850 152.360 15.170 152.690 ;
        RECT 15.330 152.660 16.360 153.190 ;
        RECT 17.090 152.690 17.820 154.040 ;
        RECT 20.380 153.390 21.320 155.220 ;
        RECT 21.570 154.760 21.830 154.790 ;
        RECT 21.570 154.470 21.850 154.760 ;
        RECT 22.010 154.670 23.010 155.220 ;
        RECT 23.880 154.790 24.610 156.140 ;
        RECT 27.100 155.560 27.450 157.390 ;
        RECT 25.330 155.290 27.450 155.560 ;
        RECT 22.010 154.500 23.010 154.510 ;
        RECT 21.570 154.450 21.830 154.470 ;
        RECT 22.000 154.290 23.010 154.500 ;
        RECT 23.150 154.460 25.180 154.790 ;
        RECT 25.340 154.760 26.370 155.290 ;
        RECT 25.355 154.730 26.355 154.760 ;
        RECT 25.355 154.500 26.355 154.520 ;
        RECT 22.000 154.200 23.150 154.290 ;
        RECT 25.330 154.200 26.370 154.500 ;
        RECT 26.530 154.460 26.850 154.790 ;
        RECT 22.000 154.060 26.370 154.200 ;
        RECT 22.000 154.040 25.380 154.060 ;
        RECT 18.690 153.120 23.010 153.390 ;
        RECT 15.345 152.630 16.345 152.660 ;
        RECT 15.345 152.400 16.345 152.420 ;
        RECT 15.330 152.100 16.370 152.400 ;
        RECT 16.520 152.360 18.550 152.690 ;
        RECT 18.690 152.570 19.690 153.120 ;
        RECT 19.870 152.660 20.130 152.690 ;
        RECT 18.690 152.400 19.690 152.410 ;
        RECT 18.690 152.190 19.700 152.400 ;
        RECT 19.850 152.370 20.130 152.660 ;
        RECT 19.870 152.350 20.130 152.370 ;
        RECT 18.550 152.100 19.700 152.190 ;
        RECT 15.330 151.960 19.700 152.100 ;
        RECT 16.320 151.940 19.700 151.960 ;
        RECT 14.250 151.090 16.370 151.360 ;
        RECT 14.250 149.260 14.600 151.090 ;
        RECT 14.850 150.260 15.170 150.590 ;
        RECT 15.330 150.560 16.360 151.090 ;
        RECT 17.090 150.590 17.820 151.940 ;
        RECT 20.380 151.290 21.320 153.120 ;
        RECT 21.570 152.660 21.830 152.690 ;
        RECT 21.570 152.370 21.850 152.660 ;
        RECT 22.010 152.570 23.010 153.120 ;
        RECT 23.880 152.690 24.610 154.040 ;
        RECT 27.100 153.460 27.450 155.290 ;
        RECT 25.330 153.190 27.450 153.460 ;
        RECT 22.010 152.400 23.010 152.410 ;
        RECT 21.570 152.350 21.830 152.370 ;
        RECT 22.000 152.190 23.010 152.400 ;
        RECT 23.150 152.360 25.180 152.690 ;
        RECT 25.340 152.660 26.370 153.190 ;
        RECT 25.355 152.630 26.355 152.660 ;
        RECT 25.355 152.400 26.355 152.420 ;
        RECT 22.000 152.100 23.150 152.190 ;
        RECT 25.330 152.100 26.370 152.400 ;
        RECT 26.530 152.360 26.850 152.690 ;
        RECT 22.000 151.960 26.370 152.100 ;
        RECT 22.000 151.940 25.380 151.960 ;
        RECT 18.690 151.020 23.010 151.290 ;
        RECT 15.345 150.530 16.345 150.560 ;
        RECT 15.345 150.300 16.345 150.320 ;
        RECT 15.330 150.000 16.370 150.300 ;
        RECT 16.520 150.260 18.550 150.590 ;
        RECT 18.690 150.470 19.690 151.020 ;
        RECT 19.870 150.560 20.130 150.590 ;
        RECT 18.690 150.300 19.690 150.310 ;
        RECT 18.690 150.090 19.700 150.300 ;
        RECT 19.850 150.270 20.130 150.560 ;
        RECT 19.870 150.250 20.130 150.270 ;
        RECT 18.550 150.000 19.700 150.090 ;
        RECT 15.330 149.860 19.700 150.000 ;
        RECT 16.320 149.840 19.700 149.860 ;
        RECT 14.250 148.990 16.370 149.260 ;
        RECT 14.250 147.160 14.600 148.990 ;
        RECT 14.850 148.160 15.170 148.490 ;
        RECT 15.330 148.460 16.360 148.990 ;
        RECT 17.090 148.490 17.820 149.840 ;
        RECT 20.380 149.190 21.320 151.020 ;
        RECT 21.570 150.560 21.830 150.590 ;
        RECT 21.570 150.270 21.850 150.560 ;
        RECT 22.010 150.470 23.010 151.020 ;
        RECT 23.880 150.590 24.610 151.940 ;
        RECT 27.100 151.360 27.450 153.190 ;
        RECT 25.330 151.090 27.450 151.360 ;
        RECT 22.010 150.300 23.010 150.310 ;
        RECT 21.570 150.250 21.830 150.270 ;
        RECT 22.000 150.090 23.010 150.300 ;
        RECT 23.150 150.260 25.180 150.590 ;
        RECT 25.340 150.560 26.370 151.090 ;
        RECT 25.355 150.530 26.355 150.560 ;
        RECT 25.355 150.300 26.355 150.320 ;
        RECT 22.000 150.000 23.150 150.090 ;
        RECT 25.330 150.000 26.370 150.300 ;
        RECT 26.530 150.260 26.850 150.590 ;
        RECT 22.000 149.860 26.370 150.000 ;
        RECT 22.000 149.840 25.380 149.860 ;
        RECT 18.690 148.920 23.010 149.190 ;
        RECT 15.345 148.430 16.345 148.460 ;
        RECT 15.345 148.200 16.345 148.220 ;
        RECT 15.330 147.900 16.370 148.200 ;
        RECT 16.520 148.160 18.550 148.490 ;
        RECT 18.690 148.370 19.690 148.920 ;
        RECT 19.870 148.460 20.130 148.490 ;
        RECT 18.690 148.200 19.690 148.210 ;
        RECT 18.690 147.990 19.700 148.200 ;
        RECT 19.850 148.170 20.130 148.460 ;
        RECT 19.870 148.150 20.130 148.170 ;
        RECT 18.550 147.900 19.700 147.990 ;
        RECT 15.330 147.760 19.700 147.900 ;
        RECT 16.320 147.740 19.700 147.760 ;
        RECT 14.250 146.890 16.370 147.160 ;
        RECT 14.250 145.060 14.600 146.890 ;
        RECT 14.850 146.060 15.170 146.390 ;
        RECT 15.330 146.360 16.360 146.890 ;
        RECT 17.090 146.390 17.820 147.740 ;
        RECT 20.380 147.090 21.320 148.920 ;
        RECT 21.570 148.460 21.830 148.490 ;
        RECT 21.570 148.170 21.850 148.460 ;
        RECT 22.010 148.370 23.010 148.920 ;
        RECT 23.880 148.490 24.610 149.840 ;
        RECT 27.100 149.260 27.450 151.090 ;
        RECT 25.330 148.990 27.450 149.260 ;
        RECT 22.010 148.200 23.010 148.210 ;
        RECT 21.570 148.150 21.830 148.170 ;
        RECT 22.000 147.990 23.010 148.200 ;
        RECT 23.150 148.160 25.180 148.490 ;
        RECT 25.340 148.460 26.370 148.990 ;
        RECT 25.355 148.430 26.355 148.460 ;
        RECT 25.355 148.200 26.355 148.220 ;
        RECT 22.000 147.900 23.150 147.990 ;
        RECT 25.330 147.900 26.370 148.200 ;
        RECT 26.530 148.160 26.850 148.490 ;
        RECT 22.000 147.760 26.370 147.900 ;
        RECT 22.000 147.740 25.380 147.760 ;
        RECT 18.690 146.820 23.010 147.090 ;
        RECT 15.345 146.330 16.345 146.360 ;
        RECT 15.345 146.100 16.345 146.120 ;
        RECT 15.330 145.800 16.370 146.100 ;
        RECT 16.520 146.060 18.550 146.390 ;
        RECT 18.690 146.270 19.690 146.820 ;
        RECT 19.870 146.360 20.130 146.390 ;
        RECT 18.690 146.100 19.690 146.110 ;
        RECT 18.690 145.890 19.700 146.100 ;
        RECT 19.850 146.070 20.130 146.360 ;
        RECT 19.870 146.050 20.130 146.070 ;
        RECT 18.550 145.800 19.700 145.890 ;
        RECT 15.330 145.660 19.700 145.800 ;
        RECT 16.320 145.640 19.700 145.660 ;
        RECT 14.250 144.790 16.370 145.060 ;
        RECT 14.250 142.960 14.600 144.790 ;
        RECT 14.850 143.960 15.170 144.290 ;
        RECT 15.330 144.260 16.360 144.790 ;
        RECT 17.090 144.290 17.820 145.640 ;
        RECT 20.380 144.990 21.320 146.820 ;
        RECT 21.570 146.360 21.830 146.390 ;
        RECT 21.570 146.070 21.850 146.360 ;
        RECT 22.010 146.270 23.010 146.820 ;
        RECT 23.880 146.390 24.610 147.740 ;
        RECT 27.100 147.160 27.450 148.990 ;
        RECT 25.330 146.890 27.450 147.160 ;
        RECT 22.010 146.100 23.010 146.110 ;
        RECT 21.570 146.050 21.830 146.070 ;
        RECT 22.000 145.890 23.010 146.100 ;
        RECT 23.150 146.060 25.180 146.390 ;
        RECT 25.340 146.360 26.370 146.890 ;
        RECT 25.355 146.330 26.355 146.360 ;
        RECT 25.355 146.100 26.355 146.120 ;
        RECT 22.000 145.800 23.150 145.890 ;
        RECT 25.330 145.800 26.370 146.100 ;
        RECT 26.530 146.060 26.850 146.390 ;
        RECT 22.000 145.660 26.370 145.800 ;
        RECT 22.000 145.640 25.380 145.660 ;
        RECT 18.690 144.720 23.010 144.990 ;
        RECT 15.345 144.230 16.345 144.260 ;
        RECT 15.345 144.000 16.345 144.020 ;
        RECT 15.330 143.700 16.370 144.000 ;
        RECT 16.520 143.960 18.550 144.290 ;
        RECT 18.690 144.170 19.690 144.720 ;
        RECT 19.870 144.260 20.130 144.290 ;
        RECT 18.690 144.000 19.690 144.010 ;
        RECT 18.690 143.790 19.700 144.000 ;
        RECT 19.850 143.970 20.130 144.260 ;
        RECT 19.870 143.950 20.130 143.970 ;
        RECT 18.550 143.700 19.700 143.790 ;
        RECT 15.330 143.560 19.700 143.700 ;
        RECT 16.320 143.540 19.700 143.560 ;
        RECT 14.250 142.690 16.370 142.960 ;
        RECT 14.250 140.860 14.600 142.690 ;
        RECT 14.850 141.860 15.170 142.190 ;
        RECT 15.330 142.160 16.360 142.690 ;
        RECT 17.090 142.190 17.820 143.540 ;
        RECT 20.380 142.890 21.320 144.720 ;
        RECT 21.570 144.260 21.830 144.290 ;
        RECT 21.570 143.970 21.850 144.260 ;
        RECT 22.010 144.170 23.010 144.720 ;
        RECT 23.880 144.290 24.610 145.640 ;
        RECT 27.100 145.060 27.450 146.890 ;
        RECT 25.330 144.790 27.450 145.060 ;
        RECT 22.010 144.000 23.010 144.010 ;
        RECT 21.570 143.950 21.830 143.970 ;
        RECT 22.000 143.790 23.010 144.000 ;
        RECT 23.150 143.960 25.180 144.290 ;
        RECT 25.340 144.260 26.370 144.790 ;
        RECT 25.355 144.230 26.355 144.260 ;
        RECT 25.355 144.000 26.355 144.020 ;
        RECT 22.000 143.700 23.150 143.790 ;
        RECT 25.330 143.700 26.370 144.000 ;
        RECT 26.530 143.960 26.850 144.290 ;
        RECT 22.000 143.560 26.370 143.700 ;
        RECT 22.000 143.540 25.380 143.560 ;
        RECT 18.690 142.620 23.010 142.890 ;
        RECT 15.345 142.130 16.345 142.160 ;
        RECT 15.345 141.900 16.345 141.920 ;
        RECT 15.330 141.600 16.370 141.900 ;
        RECT 16.520 141.860 18.550 142.190 ;
        RECT 18.690 142.070 19.690 142.620 ;
        RECT 19.870 142.160 20.130 142.190 ;
        RECT 18.690 141.900 19.690 141.910 ;
        RECT 18.690 141.690 19.700 141.900 ;
        RECT 19.850 141.870 20.130 142.160 ;
        RECT 19.870 141.850 20.130 141.870 ;
        RECT 18.550 141.600 19.700 141.690 ;
        RECT 15.330 141.460 19.700 141.600 ;
        RECT 16.320 141.440 19.700 141.460 ;
        RECT 14.250 140.590 16.370 140.860 ;
        RECT 14.250 138.760 14.600 140.590 ;
        RECT 14.850 139.760 15.170 140.090 ;
        RECT 15.330 140.060 16.360 140.590 ;
        RECT 17.090 140.090 17.820 141.440 ;
        RECT 20.380 140.790 21.320 142.620 ;
        RECT 21.570 142.160 21.830 142.190 ;
        RECT 21.570 141.870 21.850 142.160 ;
        RECT 22.010 142.070 23.010 142.620 ;
        RECT 23.880 142.190 24.610 143.540 ;
        RECT 27.100 142.960 27.450 144.790 ;
        RECT 25.330 142.690 27.450 142.960 ;
        RECT 22.010 141.900 23.010 141.910 ;
        RECT 21.570 141.850 21.830 141.870 ;
        RECT 22.000 141.690 23.010 141.900 ;
        RECT 23.150 141.860 25.180 142.190 ;
        RECT 25.340 142.160 26.370 142.690 ;
        RECT 25.355 142.130 26.355 142.160 ;
        RECT 25.355 141.900 26.355 141.920 ;
        RECT 22.000 141.600 23.150 141.690 ;
        RECT 25.330 141.600 26.370 141.900 ;
        RECT 26.530 141.860 26.850 142.190 ;
        RECT 22.000 141.460 26.370 141.600 ;
        RECT 22.000 141.440 25.380 141.460 ;
        RECT 18.690 140.520 23.010 140.790 ;
        RECT 15.345 140.030 16.345 140.060 ;
        RECT 15.345 139.800 16.345 139.820 ;
        RECT 15.330 139.500 16.370 139.800 ;
        RECT 16.520 139.760 18.550 140.090 ;
        RECT 18.690 139.970 19.690 140.520 ;
        RECT 19.870 140.060 20.130 140.090 ;
        RECT 18.690 139.800 19.690 139.810 ;
        RECT 18.690 139.590 19.700 139.800 ;
        RECT 19.850 139.770 20.130 140.060 ;
        RECT 19.870 139.750 20.130 139.770 ;
        RECT 18.550 139.500 19.700 139.590 ;
        RECT 15.330 139.360 19.700 139.500 ;
        RECT 16.320 139.340 19.700 139.360 ;
        RECT 14.250 138.490 16.370 138.760 ;
        RECT 14.250 136.660 14.600 138.490 ;
        RECT 14.850 137.660 15.170 137.990 ;
        RECT 15.330 137.960 16.360 138.490 ;
        RECT 17.090 137.990 17.820 139.340 ;
        RECT 20.380 138.690 21.320 140.520 ;
        RECT 21.570 140.060 21.830 140.090 ;
        RECT 21.570 139.770 21.850 140.060 ;
        RECT 22.010 139.970 23.010 140.520 ;
        RECT 23.880 140.090 24.610 141.440 ;
        RECT 27.100 140.860 27.450 142.690 ;
        RECT 25.330 140.590 27.450 140.860 ;
        RECT 22.010 139.800 23.010 139.810 ;
        RECT 21.570 139.750 21.830 139.770 ;
        RECT 22.000 139.590 23.010 139.800 ;
        RECT 23.150 139.760 25.180 140.090 ;
        RECT 25.340 140.060 26.370 140.590 ;
        RECT 25.355 140.030 26.355 140.060 ;
        RECT 25.355 139.800 26.355 139.820 ;
        RECT 22.000 139.500 23.150 139.590 ;
        RECT 25.330 139.500 26.370 139.800 ;
        RECT 26.530 139.760 26.850 140.090 ;
        RECT 22.000 139.360 26.370 139.500 ;
        RECT 22.000 139.340 25.380 139.360 ;
        RECT 18.690 138.420 23.010 138.690 ;
        RECT 15.345 137.930 16.345 137.960 ;
        RECT 15.345 137.700 16.345 137.720 ;
        RECT 15.330 137.400 16.370 137.700 ;
        RECT 16.520 137.660 18.550 137.990 ;
        RECT 18.690 137.870 19.690 138.420 ;
        RECT 19.870 137.960 20.130 137.990 ;
        RECT 18.690 137.700 19.690 137.710 ;
        RECT 18.690 137.490 19.700 137.700 ;
        RECT 19.850 137.670 20.130 137.960 ;
        RECT 19.870 137.650 20.130 137.670 ;
        RECT 18.550 137.400 19.700 137.490 ;
        RECT 15.330 137.260 19.700 137.400 ;
        RECT 16.320 137.240 19.700 137.260 ;
        RECT 14.250 136.390 16.370 136.660 ;
        RECT 14.250 134.560 14.600 136.390 ;
        RECT 14.850 135.560 15.170 135.890 ;
        RECT 15.330 135.860 16.360 136.390 ;
        RECT 17.090 135.890 17.820 137.240 ;
        RECT 20.380 136.590 21.320 138.420 ;
        RECT 21.570 137.960 21.830 137.990 ;
        RECT 21.570 137.670 21.850 137.960 ;
        RECT 22.010 137.870 23.010 138.420 ;
        RECT 23.880 137.990 24.610 139.340 ;
        RECT 27.100 138.760 27.450 140.590 ;
        RECT 25.330 138.490 27.450 138.760 ;
        RECT 22.010 137.700 23.010 137.710 ;
        RECT 21.570 137.650 21.830 137.670 ;
        RECT 22.000 137.490 23.010 137.700 ;
        RECT 23.150 137.660 25.180 137.990 ;
        RECT 25.340 137.960 26.370 138.490 ;
        RECT 25.355 137.930 26.355 137.960 ;
        RECT 25.355 137.700 26.355 137.720 ;
        RECT 22.000 137.400 23.150 137.490 ;
        RECT 25.330 137.400 26.370 137.700 ;
        RECT 26.530 137.660 26.850 137.990 ;
        RECT 22.000 137.260 26.370 137.400 ;
        RECT 22.000 137.240 25.380 137.260 ;
        RECT 18.690 136.320 23.010 136.590 ;
        RECT 15.345 135.830 16.345 135.860 ;
        RECT 15.345 135.600 16.345 135.620 ;
        RECT 15.330 135.300 16.370 135.600 ;
        RECT 16.520 135.560 18.550 135.890 ;
        RECT 18.690 135.770 19.690 136.320 ;
        RECT 19.870 135.860 20.130 135.890 ;
        RECT 18.690 135.600 19.690 135.610 ;
        RECT 18.690 135.390 19.700 135.600 ;
        RECT 19.850 135.570 20.130 135.860 ;
        RECT 19.870 135.550 20.130 135.570 ;
        RECT 18.550 135.300 19.700 135.390 ;
        RECT 15.330 135.160 19.700 135.300 ;
        RECT 16.320 135.140 19.700 135.160 ;
        RECT 14.250 134.290 16.370 134.560 ;
        RECT 14.250 132.460 14.600 134.290 ;
        RECT 14.850 133.460 15.170 133.790 ;
        RECT 15.330 133.760 16.360 134.290 ;
        RECT 17.090 133.790 17.820 135.140 ;
        RECT 20.380 134.490 21.320 136.320 ;
        RECT 21.570 135.860 21.830 135.890 ;
        RECT 21.570 135.570 21.850 135.860 ;
        RECT 22.010 135.770 23.010 136.320 ;
        RECT 23.880 135.890 24.610 137.240 ;
        RECT 27.100 136.660 27.450 138.490 ;
        RECT 25.330 136.390 27.450 136.660 ;
        RECT 22.010 135.600 23.010 135.610 ;
        RECT 21.570 135.550 21.830 135.570 ;
        RECT 22.000 135.390 23.010 135.600 ;
        RECT 23.150 135.560 25.180 135.890 ;
        RECT 25.340 135.860 26.370 136.390 ;
        RECT 25.355 135.830 26.355 135.860 ;
        RECT 25.355 135.600 26.355 135.620 ;
        RECT 22.000 135.300 23.150 135.390 ;
        RECT 25.330 135.300 26.370 135.600 ;
        RECT 26.530 135.560 26.850 135.890 ;
        RECT 22.000 135.160 26.370 135.300 ;
        RECT 22.000 135.140 25.380 135.160 ;
        RECT 18.690 134.220 23.010 134.490 ;
        RECT 15.345 133.730 16.345 133.760 ;
        RECT 15.345 133.500 16.345 133.520 ;
        RECT 15.330 133.200 16.370 133.500 ;
        RECT 16.520 133.460 18.550 133.790 ;
        RECT 18.690 133.670 19.690 134.220 ;
        RECT 19.870 133.760 20.130 133.790 ;
        RECT 18.690 133.500 19.690 133.510 ;
        RECT 18.690 133.290 19.700 133.500 ;
        RECT 19.850 133.470 20.130 133.760 ;
        RECT 19.870 133.450 20.130 133.470 ;
        RECT 18.550 133.200 19.700 133.290 ;
        RECT 15.330 133.060 19.700 133.200 ;
        RECT 16.320 133.040 19.700 133.060 ;
        RECT 14.250 132.190 16.370 132.460 ;
        RECT 14.250 130.360 14.600 132.190 ;
        RECT 14.850 131.360 15.170 131.690 ;
        RECT 15.330 131.660 16.360 132.190 ;
        RECT 17.090 131.690 17.820 133.040 ;
        RECT 20.380 132.390 21.320 134.220 ;
        RECT 21.570 133.760 21.830 133.790 ;
        RECT 21.570 133.470 21.850 133.760 ;
        RECT 22.010 133.670 23.010 134.220 ;
        RECT 23.880 133.790 24.610 135.140 ;
        RECT 27.100 134.560 27.450 136.390 ;
        RECT 25.330 134.290 27.450 134.560 ;
        RECT 22.010 133.500 23.010 133.510 ;
        RECT 21.570 133.450 21.830 133.470 ;
        RECT 22.000 133.290 23.010 133.500 ;
        RECT 23.150 133.460 25.180 133.790 ;
        RECT 25.340 133.760 26.370 134.290 ;
        RECT 25.355 133.730 26.355 133.760 ;
        RECT 25.355 133.500 26.355 133.520 ;
        RECT 22.000 133.200 23.150 133.290 ;
        RECT 25.330 133.200 26.370 133.500 ;
        RECT 26.530 133.460 26.850 133.790 ;
        RECT 22.000 133.060 26.370 133.200 ;
        RECT 22.000 133.040 25.380 133.060 ;
        RECT 18.690 132.120 23.010 132.390 ;
        RECT 15.345 131.630 16.345 131.660 ;
        RECT 15.345 131.400 16.345 131.420 ;
        RECT 15.330 131.100 16.370 131.400 ;
        RECT 16.520 131.360 18.550 131.690 ;
        RECT 18.690 131.570 19.690 132.120 ;
        RECT 19.870 131.660 20.130 131.690 ;
        RECT 18.690 131.400 19.690 131.410 ;
        RECT 18.690 131.190 19.700 131.400 ;
        RECT 19.850 131.370 20.130 131.660 ;
        RECT 19.870 131.350 20.130 131.370 ;
        RECT 18.550 131.100 19.700 131.190 ;
        RECT 15.330 130.960 19.700 131.100 ;
        RECT 16.320 130.940 19.700 130.960 ;
        RECT 14.250 130.090 16.370 130.360 ;
        RECT 14.250 128.260 14.600 130.090 ;
        RECT 14.850 129.260 15.170 129.590 ;
        RECT 15.330 129.560 16.360 130.090 ;
        RECT 17.090 129.590 17.820 130.940 ;
        RECT 20.380 130.290 21.320 132.120 ;
        RECT 21.570 131.660 21.830 131.690 ;
        RECT 21.570 131.370 21.850 131.660 ;
        RECT 22.010 131.570 23.010 132.120 ;
        RECT 23.880 131.690 24.610 133.040 ;
        RECT 27.100 132.460 27.450 134.290 ;
        RECT 25.330 132.190 27.450 132.460 ;
        RECT 22.010 131.400 23.010 131.410 ;
        RECT 21.570 131.350 21.830 131.370 ;
        RECT 22.000 131.190 23.010 131.400 ;
        RECT 23.150 131.360 25.180 131.690 ;
        RECT 25.340 131.660 26.370 132.190 ;
        RECT 25.355 131.630 26.355 131.660 ;
        RECT 25.355 131.400 26.355 131.420 ;
        RECT 22.000 131.100 23.150 131.190 ;
        RECT 25.330 131.100 26.370 131.400 ;
        RECT 26.530 131.360 26.850 131.690 ;
        RECT 22.000 130.960 26.370 131.100 ;
        RECT 22.000 130.940 25.380 130.960 ;
        RECT 18.690 130.020 23.010 130.290 ;
        RECT 15.345 129.530 16.345 129.560 ;
        RECT 15.345 129.300 16.345 129.320 ;
        RECT 15.330 129.000 16.370 129.300 ;
        RECT 16.520 129.260 18.550 129.590 ;
        RECT 18.690 129.470 19.690 130.020 ;
        RECT 19.870 129.560 20.130 129.590 ;
        RECT 18.690 129.300 19.690 129.310 ;
        RECT 18.690 129.090 19.700 129.300 ;
        RECT 19.850 129.270 20.130 129.560 ;
        RECT 19.870 129.250 20.130 129.270 ;
        RECT 18.550 129.000 19.700 129.090 ;
        RECT 15.330 128.860 19.700 129.000 ;
        RECT 16.320 128.840 19.700 128.860 ;
        RECT 14.250 127.990 16.370 128.260 ;
        RECT 14.250 126.160 14.600 127.990 ;
        RECT 14.850 127.160 15.170 127.490 ;
        RECT 15.330 127.460 16.360 127.990 ;
        RECT 17.090 127.490 17.820 128.840 ;
        RECT 20.380 128.190 21.320 130.020 ;
        RECT 21.570 129.560 21.830 129.590 ;
        RECT 21.570 129.270 21.850 129.560 ;
        RECT 22.010 129.470 23.010 130.020 ;
        RECT 23.880 129.590 24.610 130.940 ;
        RECT 27.100 130.360 27.450 132.190 ;
        RECT 25.330 130.090 27.450 130.360 ;
        RECT 22.010 129.300 23.010 129.310 ;
        RECT 21.570 129.250 21.830 129.270 ;
        RECT 22.000 129.090 23.010 129.300 ;
        RECT 23.150 129.260 25.180 129.590 ;
        RECT 25.340 129.560 26.370 130.090 ;
        RECT 25.355 129.530 26.355 129.560 ;
        RECT 25.355 129.300 26.355 129.320 ;
        RECT 22.000 129.000 23.150 129.090 ;
        RECT 25.330 129.000 26.370 129.300 ;
        RECT 26.530 129.260 26.850 129.590 ;
        RECT 22.000 128.860 26.370 129.000 ;
        RECT 22.000 128.840 25.380 128.860 ;
        RECT 18.690 127.920 23.010 128.190 ;
        RECT 15.345 127.430 16.345 127.460 ;
        RECT 15.345 127.200 16.345 127.220 ;
        RECT 15.330 126.900 16.370 127.200 ;
        RECT 16.520 127.160 18.550 127.490 ;
        RECT 18.690 127.370 19.690 127.920 ;
        RECT 19.870 127.460 20.130 127.490 ;
        RECT 18.690 127.200 19.690 127.210 ;
        RECT 18.690 126.990 19.700 127.200 ;
        RECT 19.850 127.170 20.130 127.460 ;
        RECT 19.870 127.150 20.130 127.170 ;
        RECT 18.550 126.900 19.700 126.990 ;
        RECT 15.330 126.760 19.700 126.900 ;
        RECT 16.320 126.740 19.700 126.760 ;
        RECT 14.250 125.890 16.370 126.160 ;
        RECT 14.250 124.060 14.600 125.890 ;
        RECT 14.850 125.060 15.170 125.390 ;
        RECT 15.330 125.360 16.360 125.890 ;
        RECT 17.090 125.390 17.820 126.740 ;
        RECT 20.380 126.090 21.320 127.920 ;
        RECT 21.570 127.460 21.830 127.490 ;
        RECT 21.570 127.170 21.850 127.460 ;
        RECT 22.010 127.370 23.010 127.920 ;
        RECT 23.880 127.490 24.610 128.840 ;
        RECT 27.100 128.260 27.450 130.090 ;
        RECT 25.330 127.990 27.450 128.260 ;
        RECT 22.010 127.200 23.010 127.210 ;
        RECT 21.570 127.150 21.830 127.170 ;
        RECT 22.000 126.990 23.010 127.200 ;
        RECT 23.150 127.160 25.180 127.490 ;
        RECT 25.340 127.460 26.370 127.990 ;
        RECT 25.355 127.430 26.355 127.460 ;
        RECT 25.355 127.200 26.355 127.220 ;
        RECT 22.000 126.900 23.150 126.990 ;
        RECT 25.330 126.900 26.370 127.200 ;
        RECT 26.530 127.160 26.850 127.490 ;
        RECT 22.000 126.760 26.370 126.900 ;
        RECT 22.000 126.740 25.380 126.760 ;
        RECT 18.690 125.820 23.010 126.090 ;
        RECT 15.345 125.330 16.345 125.360 ;
        RECT 15.345 125.100 16.345 125.120 ;
        RECT 15.330 124.800 16.370 125.100 ;
        RECT 16.520 125.060 18.550 125.390 ;
        RECT 18.690 125.270 19.690 125.820 ;
        RECT 19.870 125.360 20.130 125.390 ;
        RECT 18.690 125.100 19.690 125.110 ;
        RECT 18.690 124.890 19.700 125.100 ;
        RECT 19.850 125.070 20.130 125.360 ;
        RECT 19.870 125.050 20.130 125.070 ;
        RECT 18.550 124.800 19.700 124.890 ;
        RECT 15.330 124.660 19.700 124.800 ;
        RECT 16.320 124.640 19.700 124.660 ;
        RECT 14.250 123.790 16.370 124.060 ;
        RECT 14.250 121.960 14.600 123.790 ;
        RECT 14.850 122.960 15.170 123.290 ;
        RECT 15.330 123.260 16.360 123.790 ;
        RECT 17.090 123.290 17.820 124.640 ;
        RECT 20.380 123.990 21.320 125.820 ;
        RECT 21.570 125.360 21.830 125.390 ;
        RECT 21.570 125.070 21.850 125.360 ;
        RECT 22.010 125.270 23.010 125.820 ;
        RECT 23.880 125.390 24.610 126.740 ;
        RECT 27.100 126.160 27.450 127.990 ;
        RECT 25.330 125.890 27.450 126.160 ;
        RECT 22.010 125.100 23.010 125.110 ;
        RECT 21.570 125.050 21.830 125.070 ;
        RECT 22.000 124.890 23.010 125.100 ;
        RECT 23.150 125.060 25.180 125.390 ;
        RECT 25.340 125.360 26.370 125.890 ;
        RECT 25.355 125.330 26.355 125.360 ;
        RECT 25.355 125.100 26.355 125.120 ;
        RECT 22.000 124.800 23.150 124.890 ;
        RECT 25.330 124.800 26.370 125.100 ;
        RECT 26.530 125.060 26.850 125.390 ;
        RECT 22.000 124.660 26.370 124.800 ;
        RECT 22.000 124.640 25.380 124.660 ;
        RECT 18.690 123.720 23.010 123.990 ;
        RECT 15.345 123.230 16.345 123.260 ;
        RECT 15.345 123.000 16.345 123.020 ;
        RECT 15.330 122.700 16.370 123.000 ;
        RECT 16.520 122.960 18.550 123.290 ;
        RECT 18.690 123.170 19.690 123.720 ;
        RECT 19.870 123.260 20.130 123.290 ;
        RECT 18.690 123.000 19.690 123.010 ;
        RECT 18.690 122.790 19.700 123.000 ;
        RECT 19.850 122.970 20.130 123.260 ;
        RECT 19.870 122.950 20.130 122.970 ;
        RECT 18.550 122.700 19.700 122.790 ;
        RECT 15.330 122.560 19.700 122.700 ;
        RECT 16.320 122.540 19.700 122.560 ;
        RECT 14.250 121.690 16.370 121.960 ;
        RECT 14.250 119.860 14.600 121.690 ;
        RECT 14.850 120.860 15.170 121.190 ;
        RECT 15.330 121.160 16.360 121.690 ;
        RECT 17.090 121.190 17.820 122.540 ;
        RECT 20.380 121.890 21.320 123.720 ;
        RECT 21.570 123.260 21.830 123.290 ;
        RECT 21.570 122.970 21.850 123.260 ;
        RECT 22.010 123.170 23.010 123.720 ;
        RECT 23.880 123.290 24.610 124.640 ;
        RECT 27.100 124.060 27.450 125.890 ;
        RECT 25.330 123.790 27.450 124.060 ;
        RECT 22.010 123.000 23.010 123.010 ;
        RECT 21.570 122.950 21.830 122.970 ;
        RECT 22.000 122.790 23.010 123.000 ;
        RECT 23.150 122.960 25.180 123.290 ;
        RECT 25.340 123.260 26.370 123.790 ;
        RECT 25.355 123.230 26.355 123.260 ;
        RECT 25.355 123.000 26.355 123.020 ;
        RECT 22.000 122.700 23.150 122.790 ;
        RECT 25.330 122.700 26.370 123.000 ;
        RECT 26.530 122.960 26.850 123.290 ;
        RECT 22.000 122.560 26.370 122.700 ;
        RECT 22.000 122.540 25.380 122.560 ;
        RECT 18.690 121.620 23.010 121.890 ;
        RECT 15.345 121.130 16.345 121.160 ;
        RECT 15.345 120.900 16.345 120.920 ;
        RECT 15.330 120.600 16.370 120.900 ;
        RECT 16.520 120.860 18.550 121.190 ;
        RECT 18.690 121.070 19.690 121.620 ;
        RECT 19.870 121.160 20.130 121.190 ;
        RECT 18.690 120.900 19.690 120.910 ;
        RECT 18.690 120.690 19.700 120.900 ;
        RECT 19.850 120.870 20.130 121.160 ;
        RECT 19.870 120.850 20.130 120.870 ;
        RECT 18.550 120.600 19.700 120.690 ;
        RECT 15.330 120.460 19.700 120.600 ;
        RECT 16.320 120.440 19.700 120.460 ;
        RECT 14.250 119.590 16.370 119.860 ;
        RECT 14.250 117.760 14.600 119.590 ;
        RECT 14.850 118.760 15.170 119.090 ;
        RECT 15.330 119.060 16.360 119.590 ;
        RECT 17.090 119.090 17.820 120.440 ;
        RECT 20.380 119.790 21.320 121.620 ;
        RECT 21.570 121.160 21.830 121.190 ;
        RECT 21.570 120.870 21.850 121.160 ;
        RECT 22.010 121.070 23.010 121.620 ;
        RECT 23.880 121.190 24.610 122.540 ;
        RECT 27.100 121.960 27.450 123.790 ;
        RECT 25.330 121.690 27.450 121.960 ;
        RECT 22.010 120.900 23.010 120.910 ;
        RECT 21.570 120.850 21.830 120.870 ;
        RECT 22.000 120.690 23.010 120.900 ;
        RECT 23.150 120.860 25.180 121.190 ;
        RECT 25.340 121.160 26.370 121.690 ;
        RECT 25.355 121.130 26.355 121.160 ;
        RECT 25.355 120.900 26.355 120.920 ;
        RECT 22.000 120.600 23.150 120.690 ;
        RECT 25.330 120.600 26.370 120.900 ;
        RECT 26.530 120.860 26.850 121.190 ;
        RECT 22.000 120.460 26.370 120.600 ;
        RECT 22.000 120.440 25.380 120.460 ;
        RECT 18.690 119.520 23.010 119.790 ;
        RECT 15.345 119.030 16.345 119.060 ;
        RECT 15.345 118.800 16.345 118.820 ;
        RECT 15.330 118.500 16.370 118.800 ;
        RECT 16.520 118.760 18.550 119.090 ;
        RECT 18.690 118.970 19.690 119.520 ;
        RECT 19.870 119.060 20.130 119.090 ;
        RECT 18.690 118.800 19.690 118.810 ;
        RECT 18.690 118.590 19.700 118.800 ;
        RECT 19.850 118.770 20.130 119.060 ;
        RECT 19.870 118.750 20.130 118.770 ;
        RECT 18.550 118.500 19.700 118.590 ;
        RECT 15.330 118.360 19.700 118.500 ;
        RECT 16.320 118.340 19.700 118.360 ;
        RECT 14.250 117.490 16.370 117.760 ;
        RECT 14.250 115.660 14.600 117.490 ;
        RECT 14.850 116.660 15.170 116.990 ;
        RECT 15.330 116.960 16.360 117.490 ;
        RECT 17.090 116.990 17.820 118.340 ;
        RECT 20.380 117.690 21.320 119.520 ;
        RECT 21.570 119.060 21.830 119.090 ;
        RECT 21.570 118.770 21.850 119.060 ;
        RECT 22.010 118.970 23.010 119.520 ;
        RECT 23.880 119.090 24.610 120.440 ;
        RECT 27.100 119.860 27.450 121.690 ;
        RECT 25.330 119.590 27.450 119.860 ;
        RECT 22.010 118.800 23.010 118.810 ;
        RECT 21.570 118.750 21.830 118.770 ;
        RECT 22.000 118.590 23.010 118.800 ;
        RECT 23.150 118.760 25.180 119.090 ;
        RECT 25.340 119.060 26.370 119.590 ;
        RECT 25.355 119.030 26.355 119.060 ;
        RECT 25.355 118.800 26.355 118.820 ;
        RECT 22.000 118.500 23.150 118.590 ;
        RECT 25.330 118.500 26.370 118.800 ;
        RECT 26.530 118.760 26.850 119.090 ;
        RECT 22.000 118.360 26.370 118.500 ;
        RECT 22.000 118.340 25.380 118.360 ;
        RECT 18.690 117.420 23.010 117.690 ;
        RECT 15.345 116.930 16.345 116.960 ;
        RECT 15.345 116.700 16.345 116.720 ;
        RECT 15.330 116.400 16.370 116.700 ;
        RECT 16.520 116.660 18.550 116.990 ;
        RECT 18.690 116.870 19.690 117.420 ;
        RECT 19.870 116.960 20.130 116.990 ;
        RECT 18.690 116.700 19.690 116.710 ;
        RECT 18.690 116.490 19.700 116.700 ;
        RECT 19.850 116.670 20.130 116.960 ;
        RECT 19.870 116.650 20.130 116.670 ;
        RECT 18.550 116.400 19.700 116.490 ;
        RECT 15.330 116.260 19.700 116.400 ;
        RECT 16.320 116.240 19.700 116.260 ;
        RECT 14.250 115.390 16.370 115.660 ;
        RECT 14.250 113.560 14.600 115.390 ;
        RECT 14.850 114.560 15.170 114.890 ;
        RECT 15.330 114.860 16.360 115.390 ;
        RECT 17.090 114.890 17.820 116.240 ;
        RECT 20.380 115.590 21.320 117.420 ;
        RECT 21.570 116.960 21.830 116.990 ;
        RECT 21.570 116.670 21.850 116.960 ;
        RECT 22.010 116.870 23.010 117.420 ;
        RECT 23.880 116.990 24.610 118.340 ;
        RECT 27.100 117.760 27.450 119.590 ;
        RECT 25.330 117.490 27.450 117.760 ;
        RECT 22.010 116.700 23.010 116.710 ;
        RECT 21.570 116.650 21.830 116.670 ;
        RECT 22.000 116.490 23.010 116.700 ;
        RECT 23.150 116.660 25.180 116.990 ;
        RECT 25.340 116.960 26.370 117.490 ;
        RECT 25.355 116.930 26.355 116.960 ;
        RECT 25.355 116.700 26.355 116.720 ;
        RECT 22.000 116.400 23.150 116.490 ;
        RECT 25.330 116.400 26.370 116.700 ;
        RECT 26.530 116.660 26.850 116.990 ;
        RECT 22.000 116.260 26.370 116.400 ;
        RECT 22.000 116.240 25.380 116.260 ;
        RECT 18.690 115.320 23.010 115.590 ;
        RECT 15.345 114.830 16.345 114.860 ;
        RECT 15.345 114.600 16.345 114.620 ;
        RECT 15.330 114.300 16.370 114.600 ;
        RECT 16.520 114.560 18.550 114.890 ;
        RECT 18.690 114.770 19.690 115.320 ;
        RECT 19.870 114.860 20.130 114.890 ;
        RECT 18.690 114.600 19.690 114.610 ;
        RECT 18.690 114.390 19.700 114.600 ;
        RECT 19.850 114.570 20.130 114.860 ;
        RECT 19.870 114.550 20.130 114.570 ;
        RECT 18.550 114.300 19.700 114.390 ;
        RECT 15.330 114.160 19.700 114.300 ;
        RECT 16.320 114.140 19.700 114.160 ;
        RECT 14.250 113.290 16.370 113.560 ;
        RECT 14.250 111.460 14.600 113.290 ;
        RECT 14.850 112.460 15.170 112.790 ;
        RECT 15.330 112.760 16.360 113.290 ;
        RECT 17.090 112.790 17.820 114.140 ;
        RECT 20.380 113.490 21.320 115.320 ;
        RECT 21.570 114.860 21.830 114.890 ;
        RECT 21.570 114.570 21.850 114.860 ;
        RECT 22.010 114.770 23.010 115.320 ;
        RECT 23.880 114.890 24.610 116.240 ;
        RECT 27.100 115.660 27.450 117.490 ;
        RECT 25.330 115.390 27.450 115.660 ;
        RECT 22.010 114.600 23.010 114.610 ;
        RECT 21.570 114.550 21.830 114.570 ;
        RECT 22.000 114.390 23.010 114.600 ;
        RECT 23.150 114.560 25.180 114.890 ;
        RECT 25.340 114.860 26.370 115.390 ;
        RECT 25.355 114.830 26.355 114.860 ;
        RECT 25.355 114.600 26.355 114.620 ;
        RECT 22.000 114.300 23.150 114.390 ;
        RECT 25.330 114.300 26.370 114.600 ;
        RECT 26.530 114.560 26.850 114.890 ;
        RECT 22.000 114.160 26.370 114.300 ;
        RECT 22.000 114.140 25.380 114.160 ;
        RECT 18.690 113.220 23.010 113.490 ;
        RECT 15.345 112.730 16.345 112.760 ;
        RECT 15.345 112.500 16.345 112.520 ;
        RECT 15.330 112.200 16.370 112.500 ;
        RECT 16.520 112.460 18.550 112.790 ;
        RECT 18.690 112.670 19.690 113.220 ;
        RECT 19.870 112.760 20.130 112.790 ;
        RECT 18.690 112.500 19.690 112.510 ;
        RECT 18.690 112.290 19.700 112.500 ;
        RECT 19.850 112.470 20.130 112.760 ;
        RECT 19.870 112.450 20.130 112.470 ;
        RECT 18.550 112.200 19.700 112.290 ;
        RECT 15.330 112.060 19.700 112.200 ;
        RECT 16.320 112.040 19.700 112.060 ;
        RECT 14.250 111.190 16.370 111.460 ;
        RECT 14.250 109.360 14.600 111.190 ;
        RECT 14.850 110.360 15.170 110.690 ;
        RECT 15.330 110.660 16.360 111.190 ;
        RECT 17.090 110.690 17.820 112.040 ;
        RECT 20.380 111.390 21.320 113.220 ;
        RECT 21.570 112.760 21.830 112.790 ;
        RECT 21.570 112.470 21.850 112.760 ;
        RECT 22.010 112.670 23.010 113.220 ;
        RECT 23.880 112.790 24.610 114.140 ;
        RECT 27.100 113.560 27.450 115.390 ;
        RECT 25.330 113.290 27.450 113.560 ;
        RECT 22.010 112.500 23.010 112.510 ;
        RECT 21.570 112.450 21.830 112.470 ;
        RECT 22.000 112.290 23.010 112.500 ;
        RECT 23.150 112.460 25.180 112.790 ;
        RECT 25.340 112.760 26.370 113.290 ;
        RECT 25.355 112.730 26.355 112.760 ;
        RECT 25.355 112.500 26.355 112.520 ;
        RECT 22.000 112.200 23.150 112.290 ;
        RECT 25.330 112.200 26.370 112.500 ;
        RECT 26.530 112.460 26.850 112.790 ;
        RECT 22.000 112.060 26.370 112.200 ;
        RECT 22.000 112.040 25.380 112.060 ;
        RECT 18.690 111.120 23.010 111.390 ;
        RECT 15.345 110.630 16.345 110.660 ;
        RECT 15.345 110.400 16.345 110.420 ;
        RECT 15.330 110.100 16.370 110.400 ;
        RECT 16.520 110.360 18.550 110.690 ;
        RECT 18.690 110.570 19.690 111.120 ;
        RECT 19.870 110.660 20.130 110.690 ;
        RECT 18.690 110.400 19.690 110.410 ;
        RECT 18.690 110.190 19.700 110.400 ;
        RECT 19.850 110.370 20.130 110.660 ;
        RECT 19.870 110.350 20.130 110.370 ;
        RECT 18.550 110.100 19.700 110.190 ;
        RECT 15.330 109.960 19.700 110.100 ;
        RECT 16.320 109.940 19.700 109.960 ;
        RECT 14.250 109.090 16.370 109.360 ;
        RECT 14.250 107.260 14.600 109.090 ;
        RECT 14.850 108.260 15.170 108.590 ;
        RECT 15.330 108.560 16.360 109.090 ;
        RECT 17.090 108.590 17.820 109.940 ;
        RECT 20.380 109.290 21.320 111.120 ;
        RECT 21.570 110.660 21.830 110.690 ;
        RECT 21.570 110.370 21.850 110.660 ;
        RECT 22.010 110.570 23.010 111.120 ;
        RECT 23.880 110.690 24.610 112.040 ;
        RECT 27.100 111.460 27.450 113.290 ;
        RECT 25.330 111.190 27.450 111.460 ;
        RECT 22.010 110.400 23.010 110.410 ;
        RECT 21.570 110.350 21.830 110.370 ;
        RECT 22.000 110.190 23.010 110.400 ;
        RECT 23.150 110.360 25.180 110.690 ;
        RECT 25.340 110.660 26.370 111.190 ;
        RECT 25.355 110.630 26.355 110.660 ;
        RECT 25.355 110.400 26.355 110.420 ;
        RECT 22.000 110.100 23.150 110.190 ;
        RECT 25.330 110.100 26.370 110.400 ;
        RECT 26.530 110.360 26.850 110.690 ;
        RECT 22.000 109.960 26.370 110.100 ;
        RECT 22.000 109.940 25.380 109.960 ;
        RECT 18.690 109.020 23.010 109.290 ;
        RECT 15.345 108.530 16.345 108.560 ;
        RECT 15.345 108.300 16.345 108.320 ;
        RECT 15.330 108.000 16.370 108.300 ;
        RECT 16.520 108.260 18.550 108.590 ;
        RECT 18.690 108.470 19.690 109.020 ;
        RECT 19.870 108.560 20.130 108.590 ;
        RECT 18.690 108.300 19.690 108.310 ;
        RECT 18.690 108.090 19.700 108.300 ;
        RECT 19.850 108.270 20.130 108.560 ;
        RECT 19.870 108.250 20.130 108.270 ;
        RECT 18.550 108.000 19.700 108.090 ;
        RECT 15.330 107.860 19.700 108.000 ;
        RECT 16.320 107.840 19.700 107.860 ;
        RECT 14.250 106.990 16.370 107.260 ;
        RECT 14.250 105.160 14.600 106.990 ;
        RECT 14.850 106.160 15.170 106.490 ;
        RECT 15.330 106.460 16.360 106.990 ;
        RECT 17.090 106.490 17.820 107.840 ;
        RECT 20.380 107.190 21.320 109.020 ;
        RECT 21.570 108.560 21.830 108.590 ;
        RECT 21.570 108.270 21.850 108.560 ;
        RECT 22.010 108.470 23.010 109.020 ;
        RECT 23.880 108.590 24.610 109.940 ;
        RECT 27.100 109.360 27.450 111.190 ;
        RECT 25.330 109.090 27.450 109.360 ;
        RECT 22.010 108.300 23.010 108.310 ;
        RECT 21.570 108.250 21.830 108.270 ;
        RECT 22.000 108.090 23.010 108.300 ;
        RECT 23.150 108.260 25.180 108.590 ;
        RECT 25.340 108.560 26.370 109.090 ;
        RECT 25.355 108.530 26.355 108.560 ;
        RECT 25.355 108.300 26.355 108.320 ;
        RECT 22.000 108.000 23.150 108.090 ;
        RECT 25.330 108.000 26.370 108.300 ;
        RECT 26.530 108.260 26.850 108.590 ;
        RECT 22.000 107.860 26.370 108.000 ;
        RECT 22.000 107.840 25.380 107.860 ;
        RECT 18.690 106.920 23.010 107.190 ;
        RECT 15.345 106.430 16.345 106.460 ;
        RECT 15.345 106.200 16.345 106.220 ;
        RECT 15.330 105.900 16.370 106.200 ;
        RECT 16.520 106.160 18.550 106.490 ;
        RECT 18.690 106.370 19.690 106.920 ;
        RECT 19.870 106.460 20.130 106.490 ;
        RECT 18.690 106.200 19.690 106.210 ;
        RECT 18.690 105.990 19.700 106.200 ;
        RECT 19.850 106.170 20.130 106.460 ;
        RECT 19.870 106.150 20.130 106.170 ;
        RECT 18.550 105.900 19.700 105.990 ;
        RECT 15.330 105.760 19.700 105.900 ;
        RECT 16.320 105.740 19.700 105.760 ;
        RECT 14.250 104.890 16.370 105.160 ;
        RECT 14.250 103.060 14.600 104.890 ;
        RECT 14.850 104.060 15.170 104.390 ;
        RECT 15.330 104.360 16.360 104.890 ;
        RECT 17.090 104.390 17.820 105.740 ;
        RECT 20.380 105.090 21.320 106.920 ;
        RECT 21.570 106.460 21.830 106.490 ;
        RECT 21.570 106.170 21.850 106.460 ;
        RECT 22.010 106.370 23.010 106.920 ;
        RECT 23.880 106.490 24.610 107.840 ;
        RECT 27.100 107.260 27.450 109.090 ;
        RECT 25.330 106.990 27.450 107.260 ;
        RECT 22.010 106.200 23.010 106.210 ;
        RECT 21.570 106.150 21.830 106.170 ;
        RECT 22.000 105.990 23.010 106.200 ;
        RECT 23.150 106.160 25.180 106.490 ;
        RECT 25.340 106.460 26.370 106.990 ;
        RECT 25.355 106.430 26.355 106.460 ;
        RECT 25.355 106.200 26.355 106.220 ;
        RECT 22.000 105.900 23.150 105.990 ;
        RECT 25.330 105.900 26.370 106.200 ;
        RECT 26.530 106.160 26.850 106.490 ;
        RECT 22.000 105.760 26.370 105.900 ;
        RECT 22.000 105.740 25.380 105.760 ;
        RECT 18.690 104.820 23.010 105.090 ;
        RECT 15.345 104.330 16.345 104.360 ;
        RECT 15.345 104.100 16.345 104.120 ;
        RECT 15.330 103.800 16.370 104.100 ;
        RECT 16.520 104.060 18.550 104.390 ;
        RECT 18.690 104.270 19.690 104.820 ;
        RECT 19.870 104.360 20.130 104.390 ;
        RECT 18.690 104.100 19.690 104.110 ;
        RECT 18.690 103.890 19.700 104.100 ;
        RECT 19.850 104.070 20.130 104.360 ;
        RECT 19.870 104.050 20.130 104.070 ;
        RECT 18.550 103.800 19.700 103.890 ;
        RECT 15.330 103.660 19.700 103.800 ;
        RECT 16.320 103.640 19.700 103.660 ;
        RECT 14.250 102.790 16.370 103.060 ;
        RECT 14.250 100.960 14.600 102.790 ;
        RECT 14.850 101.960 15.170 102.290 ;
        RECT 15.330 102.260 16.360 102.790 ;
        RECT 17.090 102.290 17.820 103.640 ;
        RECT 20.380 102.990 21.320 104.820 ;
        RECT 21.570 104.360 21.830 104.390 ;
        RECT 21.570 104.070 21.850 104.360 ;
        RECT 22.010 104.270 23.010 104.820 ;
        RECT 23.880 104.390 24.610 105.740 ;
        RECT 27.100 105.160 27.450 106.990 ;
        RECT 25.330 104.890 27.450 105.160 ;
        RECT 22.010 104.100 23.010 104.110 ;
        RECT 21.570 104.050 21.830 104.070 ;
        RECT 22.000 103.890 23.010 104.100 ;
        RECT 23.150 104.060 25.180 104.390 ;
        RECT 25.340 104.360 26.370 104.890 ;
        RECT 25.355 104.330 26.355 104.360 ;
        RECT 25.355 104.100 26.355 104.120 ;
        RECT 22.000 103.800 23.150 103.890 ;
        RECT 25.330 103.800 26.370 104.100 ;
        RECT 26.530 104.060 26.850 104.390 ;
        RECT 22.000 103.660 26.370 103.800 ;
        RECT 22.000 103.640 25.380 103.660 ;
        RECT 18.690 102.720 23.010 102.990 ;
        RECT 15.345 102.230 16.345 102.260 ;
        RECT 15.345 102.000 16.345 102.020 ;
        RECT 15.330 101.700 16.370 102.000 ;
        RECT 16.520 101.960 18.550 102.290 ;
        RECT 18.690 102.170 19.690 102.720 ;
        RECT 19.870 102.260 20.130 102.290 ;
        RECT 18.690 102.000 19.690 102.010 ;
        RECT 18.690 101.790 19.700 102.000 ;
        RECT 19.850 101.970 20.130 102.260 ;
        RECT 19.870 101.950 20.130 101.970 ;
        RECT 18.550 101.700 19.700 101.790 ;
        RECT 15.330 101.560 19.700 101.700 ;
        RECT 16.320 101.540 19.700 101.560 ;
        RECT 14.250 100.690 16.370 100.960 ;
        RECT 14.250 98.860 14.600 100.690 ;
        RECT 14.850 99.860 15.170 100.190 ;
        RECT 15.330 100.160 16.360 100.690 ;
        RECT 17.090 100.190 17.820 101.540 ;
        RECT 20.380 100.890 21.320 102.720 ;
        RECT 21.570 102.260 21.830 102.290 ;
        RECT 21.570 101.970 21.850 102.260 ;
        RECT 22.010 102.170 23.010 102.720 ;
        RECT 23.880 102.290 24.610 103.640 ;
        RECT 27.100 103.060 27.450 104.890 ;
        RECT 25.330 102.790 27.450 103.060 ;
        RECT 22.010 102.000 23.010 102.010 ;
        RECT 21.570 101.950 21.830 101.970 ;
        RECT 22.000 101.790 23.010 102.000 ;
        RECT 23.150 101.960 25.180 102.290 ;
        RECT 25.340 102.260 26.370 102.790 ;
        RECT 25.355 102.230 26.355 102.260 ;
        RECT 25.355 102.000 26.355 102.020 ;
        RECT 22.000 101.700 23.150 101.790 ;
        RECT 25.330 101.700 26.370 102.000 ;
        RECT 26.530 101.960 26.850 102.290 ;
        RECT 22.000 101.560 26.370 101.700 ;
        RECT 22.000 101.540 25.380 101.560 ;
        RECT 18.690 100.620 23.010 100.890 ;
        RECT 15.345 100.130 16.345 100.160 ;
        RECT 15.345 99.900 16.345 99.920 ;
        RECT 15.330 99.600 16.370 99.900 ;
        RECT 16.520 99.860 18.550 100.190 ;
        RECT 18.690 100.070 19.690 100.620 ;
        RECT 19.870 100.160 20.130 100.190 ;
        RECT 18.690 99.900 19.690 99.910 ;
        RECT 18.690 99.690 19.700 99.900 ;
        RECT 19.850 99.870 20.130 100.160 ;
        RECT 19.870 99.850 20.130 99.870 ;
        RECT 18.550 99.600 19.700 99.690 ;
        RECT 15.330 99.460 19.700 99.600 ;
        RECT 16.320 99.440 19.700 99.460 ;
        RECT 14.250 98.590 16.370 98.860 ;
        RECT 14.250 96.760 14.600 98.590 ;
        RECT 14.850 97.760 15.170 98.090 ;
        RECT 15.330 98.060 16.360 98.590 ;
        RECT 17.090 98.090 17.820 99.440 ;
        RECT 20.380 98.790 21.320 100.620 ;
        RECT 21.570 100.160 21.830 100.190 ;
        RECT 21.570 99.870 21.850 100.160 ;
        RECT 22.010 100.070 23.010 100.620 ;
        RECT 23.880 100.190 24.610 101.540 ;
        RECT 27.100 100.960 27.450 102.790 ;
        RECT 25.330 100.690 27.450 100.960 ;
        RECT 22.010 99.900 23.010 99.910 ;
        RECT 21.570 99.850 21.830 99.870 ;
        RECT 22.000 99.690 23.010 99.900 ;
        RECT 23.150 99.860 25.180 100.190 ;
        RECT 25.340 100.160 26.370 100.690 ;
        RECT 25.355 100.130 26.355 100.160 ;
        RECT 25.355 99.900 26.355 99.920 ;
        RECT 22.000 99.600 23.150 99.690 ;
        RECT 25.330 99.600 26.370 99.900 ;
        RECT 26.530 99.860 26.850 100.190 ;
        RECT 22.000 99.460 26.370 99.600 ;
        RECT 22.000 99.440 25.380 99.460 ;
        RECT 18.690 98.520 23.010 98.790 ;
        RECT 15.345 98.030 16.345 98.060 ;
        RECT 15.345 97.800 16.345 97.820 ;
        RECT 15.330 97.500 16.370 97.800 ;
        RECT 16.520 97.760 18.550 98.090 ;
        RECT 18.690 97.970 19.690 98.520 ;
        RECT 19.870 98.060 20.130 98.090 ;
        RECT 18.690 97.800 19.690 97.810 ;
        RECT 18.690 97.590 19.700 97.800 ;
        RECT 19.850 97.770 20.130 98.060 ;
        RECT 19.870 97.750 20.130 97.770 ;
        RECT 18.550 97.500 19.700 97.590 ;
        RECT 15.330 97.360 19.700 97.500 ;
        RECT 16.320 97.340 19.700 97.360 ;
        RECT 14.250 96.490 16.370 96.760 ;
        RECT 14.250 94.660 14.600 96.490 ;
        RECT 14.850 95.660 15.170 95.990 ;
        RECT 15.330 95.960 16.360 96.490 ;
        RECT 17.090 95.990 17.820 97.340 ;
        RECT 20.380 96.690 21.320 98.520 ;
        RECT 21.570 98.060 21.830 98.090 ;
        RECT 21.570 97.770 21.850 98.060 ;
        RECT 22.010 97.970 23.010 98.520 ;
        RECT 23.880 98.090 24.610 99.440 ;
        RECT 27.100 98.860 27.450 100.690 ;
        RECT 25.330 98.590 27.450 98.860 ;
        RECT 22.010 97.800 23.010 97.810 ;
        RECT 21.570 97.750 21.830 97.770 ;
        RECT 22.000 97.590 23.010 97.800 ;
        RECT 23.150 97.760 25.180 98.090 ;
        RECT 25.340 98.060 26.370 98.590 ;
        RECT 25.355 98.030 26.355 98.060 ;
        RECT 25.355 97.800 26.355 97.820 ;
        RECT 22.000 97.500 23.150 97.590 ;
        RECT 25.330 97.500 26.370 97.800 ;
        RECT 26.530 97.760 26.850 98.090 ;
        RECT 22.000 97.360 26.370 97.500 ;
        RECT 22.000 97.340 25.380 97.360 ;
        RECT 18.690 96.420 23.010 96.690 ;
        RECT 15.345 95.930 16.345 95.960 ;
        RECT 15.345 95.700 16.345 95.720 ;
        RECT 15.330 95.400 16.370 95.700 ;
        RECT 16.520 95.660 18.550 95.990 ;
        RECT 18.690 95.870 19.690 96.420 ;
        RECT 19.870 95.960 20.130 95.990 ;
        RECT 18.690 95.700 19.690 95.710 ;
        RECT 18.690 95.490 19.700 95.700 ;
        RECT 19.850 95.670 20.130 95.960 ;
        RECT 19.870 95.650 20.130 95.670 ;
        RECT 18.550 95.400 19.700 95.490 ;
        RECT 15.330 95.260 19.700 95.400 ;
        RECT 16.320 95.240 19.700 95.260 ;
        RECT 14.250 94.390 16.370 94.660 ;
        RECT 14.250 92.560 14.600 94.390 ;
        RECT 14.850 93.560 15.170 93.890 ;
        RECT 15.330 93.860 16.360 94.390 ;
        RECT 17.090 93.890 17.820 95.240 ;
        RECT 20.380 94.590 21.320 96.420 ;
        RECT 21.570 95.960 21.830 95.990 ;
        RECT 21.570 95.670 21.850 95.960 ;
        RECT 22.010 95.870 23.010 96.420 ;
        RECT 23.880 95.990 24.610 97.340 ;
        RECT 27.100 96.760 27.450 98.590 ;
        RECT 25.330 96.490 27.450 96.760 ;
        RECT 22.010 95.700 23.010 95.710 ;
        RECT 21.570 95.650 21.830 95.670 ;
        RECT 22.000 95.490 23.010 95.700 ;
        RECT 23.150 95.660 25.180 95.990 ;
        RECT 25.340 95.960 26.370 96.490 ;
        RECT 25.355 95.930 26.355 95.960 ;
        RECT 25.355 95.700 26.355 95.720 ;
        RECT 22.000 95.400 23.150 95.490 ;
        RECT 25.330 95.400 26.370 95.700 ;
        RECT 26.530 95.660 26.850 95.990 ;
        RECT 22.000 95.260 26.370 95.400 ;
        RECT 22.000 95.240 25.380 95.260 ;
        RECT 18.690 94.320 23.010 94.590 ;
        RECT 15.345 93.830 16.345 93.860 ;
        RECT 15.345 93.600 16.345 93.620 ;
        RECT 15.330 93.300 16.370 93.600 ;
        RECT 16.520 93.560 18.550 93.890 ;
        RECT 18.690 93.770 19.690 94.320 ;
        RECT 19.870 93.860 20.130 93.890 ;
        RECT 18.690 93.600 19.690 93.610 ;
        RECT 18.690 93.390 19.700 93.600 ;
        RECT 19.850 93.570 20.130 93.860 ;
        RECT 19.870 93.550 20.130 93.570 ;
        RECT 18.550 93.300 19.700 93.390 ;
        RECT 15.330 93.160 19.700 93.300 ;
        RECT 16.320 93.140 19.700 93.160 ;
        RECT 14.250 92.290 16.370 92.560 ;
        RECT 14.250 90.460 14.600 92.290 ;
        RECT 14.850 91.460 15.170 91.790 ;
        RECT 15.330 91.760 16.360 92.290 ;
        RECT 17.090 91.790 17.820 93.140 ;
        RECT 20.380 92.490 21.320 94.320 ;
        RECT 21.570 93.860 21.830 93.890 ;
        RECT 21.570 93.570 21.850 93.860 ;
        RECT 22.010 93.770 23.010 94.320 ;
        RECT 23.880 93.890 24.610 95.240 ;
        RECT 27.100 94.660 27.450 96.490 ;
        RECT 25.330 94.390 27.450 94.660 ;
        RECT 22.010 93.600 23.010 93.610 ;
        RECT 21.570 93.550 21.830 93.570 ;
        RECT 22.000 93.390 23.010 93.600 ;
        RECT 23.150 93.560 25.180 93.890 ;
        RECT 25.340 93.860 26.370 94.390 ;
        RECT 25.355 93.830 26.355 93.860 ;
        RECT 25.355 93.600 26.355 93.620 ;
        RECT 22.000 93.300 23.150 93.390 ;
        RECT 25.330 93.300 26.370 93.600 ;
        RECT 26.530 93.560 26.850 93.890 ;
        RECT 22.000 93.160 26.370 93.300 ;
        RECT 22.000 93.140 25.380 93.160 ;
        RECT 18.690 92.220 23.010 92.490 ;
        RECT 15.345 91.730 16.345 91.760 ;
        RECT 15.345 91.500 16.345 91.520 ;
        RECT 15.330 91.200 16.370 91.500 ;
        RECT 16.520 91.460 18.550 91.790 ;
        RECT 18.690 91.670 19.690 92.220 ;
        RECT 19.870 91.760 20.130 91.790 ;
        RECT 18.690 91.500 19.690 91.510 ;
        RECT 18.690 91.290 19.700 91.500 ;
        RECT 19.850 91.470 20.130 91.760 ;
        RECT 19.870 91.450 20.130 91.470 ;
        RECT 18.550 91.200 19.700 91.290 ;
        RECT 15.330 91.060 19.700 91.200 ;
        RECT 16.320 91.040 19.700 91.060 ;
        RECT 14.250 90.190 16.370 90.460 ;
        RECT 14.250 88.360 14.600 90.190 ;
        RECT 14.850 89.360 15.170 89.690 ;
        RECT 15.330 89.660 16.360 90.190 ;
        RECT 17.090 89.690 17.820 91.040 ;
        RECT 20.380 90.390 21.320 92.220 ;
        RECT 21.570 91.760 21.830 91.790 ;
        RECT 21.570 91.470 21.850 91.760 ;
        RECT 22.010 91.670 23.010 92.220 ;
        RECT 23.880 91.790 24.610 93.140 ;
        RECT 27.100 92.560 27.450 94.390 ;
        RECT 25.330 92.290 27.450 92.560 ;
        RECT 22.010 91.500 23.010 91.510 ;
        RECT 21.570 91.450 21.830 91.470 ;
        RECT 22.000 91.290 23.010 91.500 ;
        RECT 23.150 91.460 25.180 91.790 ;
        RECT 25.340 91.760 26.370 92.290 ;
        RECT 25.355 91.730 26.355 91.760 ;
        RECT 25.355 91.500 26.355 91.520 ;
        RECT 22.000 91.200 23.150 91.290 ;
        RECT 25.330 91.200 26.370 91.500 ;
        RECT 26.530 91.460 26.850 91.790 ;
        RECT 22.000 91.060 26.370 91.200 ;
        RECT 22.000 91.040 25.380 91.060 ;
        RECT 18.690 90.120 23.010 90.390 ;
        RECT 15.345 89.630 16.345 89.660 ;
        RECT 15.345 89.400 16.345 89.420 ;
        RECT 15.330 89.100 16.370 89.400 ;
        RECT 16.520 89.360 18.550 89.690 ;
        RECT 18.690 89.570 19.690 90.120 ;
        RECT 19.870 89.660 20.130 89.690 ;
        RECT 18.690 89.400 19.690 89.410 ;
        RECT 18.690 89.190 19.700 89.400 ;
        RECT 19.850 89.370 20.130 89.660 ;
        RECT 19.870 89.350 20.130 89.370 ;
        RECT 18.550 89.100 19.700 89.190 ;
        RECT 15.330 88.960 19.700 89.100 ;
        RECT 16.320 88.940 19.700 88.960 ;
        RECT 14.250 88.090 16.370 88.360 ;
        RECT 14.250 86.260 14.600 88.090 ;
        RECT 14.850 87.260 15.170 87.590 ;
        RECT 15.330 87.560 16.360 88.090 ;
        RECT 17.090 87.590 17.820 88.940 ;
        RECT 20.380 88.290 21.320 90.120 ;
        RECT 21.570 89.660 21.830 89.690 ;
        RECT 21.570 89.370 21.850 89.660 ;
        RECT 22.010 89.570 23.010 90.120 ;
        RECT 23.880 89.690 24.610 91.040 ;
        RECT 27.100 90.460 27.450 92.290 ;
        RECT 25.330 90.190 27.450 90.460 ;
        RECT 22.010 89.400 23.010 89.410 ;
        RECT 21.570 89.350 21.830 89.370 ;
        RECT 22.000 89.190 23.010 89.400 ;
        RECT 23.150 89.360 25.180 89.690 ;
        RECT 25.340 89.660 26.370 90.190 ;
        RECT 25.355 89.630 26.355 89.660 ;
        RECT 25.355 89.400 26.355 89.420 ;
        RECT 22.000 89.100 23.150 89.190 ;
        RECT 25.330 89.100 26.370 89.400 ;
        RECT 26.530 89.360 26.850 89.690 ;
        RECT 22.000 88.960 26.370 89.100 ;
        RECT 22.000 88.940 25.380 88.960 ;
        RECT 18.690 88.020 23.010 88.290 ;
        RECT 15.345 87.530 16.345 87.560 ;
        RECT 15.345 87.300 16.345 87.320 ;
        RECT 15.330 87.000 16.370 87.300 ;
        RECT 16.520 87.260 18.550 87.590 ;
        RECT 18.690 87.470 19.690 88.020 ;
        RECT 19.870 87.560 20.130 87.590 ;
        RECT 18.690 87.300 19.690 87.310 ;
        RECT 18.690 87.090 19.700 87.300 ;
        RECT 19.850 87.270 20.130 87.560 ;
        RECT 19.870 87.250 20.130 87.270 ;
        RECT 18.550 87.000 19.700 87.090 ;
        RECT 15.330 86.860 19.700 87.000 ;
        RECT 16.320 86.840 19.700 86.860 ;
        RECT 14.250 85.990 16.370 86.260 ;
        RECT 14.250 84.160 14.600 85.990 ;
        RECT 14.850 85.160 15.170 85.490 ;
        RECT 15.330 85.460 16.360 85.990 ;
        RECT 17.090 85.490 17.820 86.840 ;
        RECT 20.380 86.190 21.320 88.020 ;
        RECT 21.570 87.560 21.830 87.590 ;
        RECT 21.570 87.270 21.850 87.560 ;
        RECT 22.010 87.470 23.010 88.020 ;
        RECT 23.880 87.590 24.610 88.940 ;
        RECT 27.100 88.360 27.450 90.190 ;
        RECT 25.330 88.090 27.450 88.360 ;
        RECT 22.010 87.300 23.010 87.310 ;
        RECT 21.570 87.250 21.830 87.270 ;
        RECT 22.000 87.090 23.010 87.300 ;
        RECT 23.150 87.260 25.180 87.590 ;
        RECT 25.340 87.560 26.370 88.090 ;
        RECT 25.355 87.530 26.355 87.560 ;
        RECT 25.355 87.300 26.355 87.320 ;
        RECT 22.000 87.000 23.150 87.090 ;
        RECT 25.330 87.000 26.370 87.300 ;
        RECT 26.530 87.260 26.850 87.590 ;
        RECT 22.000 86.860 26.370 87.000 ;
        RECT 22.000 86.840 25.380 86.860 ;
        RECT 18.690 85.920 23.010 86.190 ;
        RECT 15.345 85.430 16.345 85.460 ;
        RECT 15.345 85.200 16.345 85.220 ;
        RECT 15.330 84.900 16.370 85.200 ;
        RECT 16.520 85.160 18.550 85.490 ;
        RECT 18.690 85.370 19.690 85.920 ;
        RECT 19.870 85.460 20.130 85.490 ;
        RECT 18.690 85.200 19.690 85.210 ;
        RECT 18.690 84.990 19.700 85.200 ;
        RECT 19.850 85.170 20.130 85.460 ;
        RECT 19.870 85.150 20.130 85.170 ;
        RECT 18.550 84.900 19.700 84.990 ;
        RECT 15.330 84.760 19.700 84.900 ;
        RECT 16.320 84.740 19.700 84.760 ;
        RECT 14.250 83.890 16.370 84.160 ;
        RECT 14.250 82.060 14.600 83.890 ;
        RECT 14.850 83.060 15.170 83.390 ;
        RECT 15.330 83.360 16.360 83.890 ;
        RECT 17.090 83.390 17.820 84.740 ;
        RECT 20.380 84.090 21.320 85.920 ;
        RECT 21.570 85.460 21.830 85.490 ;
        RECT 21.570 85.170 21.850 85.460 ;
        RECT 22.010 85.370 23.010 85.920 ;
        RECT 23.880 85.490 24.610 86.840 ;
        RECT 27.100 86.260 27.450 88.090 ;
        RECT 25.330 85.990 27.450 86.260 ;
        RECT 22.010 85.200 23.010 85.210 ;
        RECT 21.570 85.150 21.830 85.170 ;
        RECT 22.000 84.990 23.010 85.200 ;
        RECT 23.150 85.160 25.180 85.490 ;
        RECT 25.340 85.460 26.370 85.990 ;
        RECT 25.355 85.430 26.355 85.460 ;
        RECT 25.355 85.200 26.355 85.220 ;
        RECT 22.000 84.900 23.150 84.990 ;
        RECT 25.330 84.900 26.370 85.200 ;
        RECT 26.530 85.160 26.850 85.490 ;
        RECT 22.000 84.760 26.370 84.900 ;
        RECT 22.000 84.740 25.380 84.760 ;
        RECT 18.690 83.820 23.010 84.090 ;
        RECT 15.345 83.330 16.345 83.360 ;
        RECT 15.345 83.100 16.345 83.120 ;
        RECT 15.330 82.800 16.370 83.100 ;
        RECT 16.520 83.060 18.550 83.390 ;
        RECT 18.690 83.270 19.690 83.820 ;
        RECT 19.870 83.360 20.130 83.390 ;
        RECT 18.690 83.100 19.690 83.110 ;
        RECT 18.690 82.890 19.700 83.100 ;
        RECT 19.850 83.070 20.130 83.360 ;
        RECT 19.870 83.050 20.130 83.070 ;
        RECT 18.550 82.800 19.700 82.890 ;
        RECT 15.330 82.660 19.700 82.800 ;
        RECT 16.320 82.640 19.700 82.660 ;
        RECT 14.250 81.790 16.370 82.060 ;
        RECT 14.250 79.960 14.600 81.790 ;
        RECT 14.850 80.960 15.170 81.290 ;
        RECT 15.330 81.260 16.360 81.790 ;
        RECT 17.090 81.290 17.820 82.640 ;
        RECT 20.380 81.990 21.320 83.820 ;
        RECT 21.570 83.360 21.830 83.390 ;
        RECT 21.570 83.070 21.850 83.360 ;
        RECT 22.010 83.270 23.010 83.820 ;
        RECT 23.880 83.390 24.610 84.740 ;
        RECT 27.100 84.160 27.450 85.990 ;
        RECT 25.330 83.890 27.450 84.160 ;
        RECT 22.010 83.100 23.010 83.110 ;
        RECT 21.570 83.050 21.830 83.070 ;
        RECT 22.000 82.890 23.010 83.100 ;
        RECT 23.150 83.060 25.180 83.390 ;
        RECT 25.340 83.360 26.370 83.890 ;
        RECT 25.355 83.330 26.355 83.360 ;
        RECT 25.355 83.100 26.355 83.120 ;
        RECT 22.000 82.800 23.150 82.890 ;
        RECT 25.330 82.800 26.370 83.100 ;
        RECT 26.530 83.060 26.850 83.390 ;
        RECT 22.000 82.660 26.370 82.800 ;
        RECT 22.000 82.640 25.380 82.660 ;
        RECT 18.690 81.720 23.010 81.990 ;
        RECT 15.345 81.230 16.345 81.260 ;
        RECT 15.345 81.000 16.345 81.020 ;
        RECT 15.330 80.700 16.370 81.000 ;
        RECT 16.520 80.960 18.550 81.290 ;
        RECT 18.690 81.170 19.690 81.720 ;
        RECT 19.870 81.260 20.130 81.290 ;
        RECT 18.690 81.000 19.690 81.010 ;
        RECT 18.690 80.790 19.700 81.000 ;
        RECT 19.850 80.970 20.130 81.260 ;
        RECT 19.870 80.950 20.130 80.970 ;
        RECT 18.550 80.700 19.700 80.790 ;
        RECT 15.330 80.560 19.700 80.700 ;
        RECT 16.320 80.540 19.700 80.560 ;
        RECT 14.250 79.690 16.370 79.960 ;
        RECT 14.250 77.860 14.600 79.690 ;
        RECT 14.850 78.860 15.170 79.190 ;
        RECT 15.330 79.160 16.360 79.690 ;
        RECT 17.090 79.190 17.820 80.540 ;
        RECT 20.380 79.890 21.320 81.720 ;
        RECT 21.570 81.260 21.830 81.290 ;
        RECT 21.570 80.970 21.850 81.260 ;
        RECT 22.010 81.170 23.010 81.720 ;
        RECT 23.880 81.290 24.610 82.640 ;
        RECT 27.100 82.060 27.450 83.890 ;
        RECT 25.330 81.790 27.450 82.060 ;
        RECT 22.010 81.000 23.010 81.010 ;
        RECT 21.570 80.950 21.830 80.970 ;
        RECT 22.000 80.790 23.010 81.000 ;
        RECT 23.150 80.960 25.180 81.290 ;
        RECT 25.340 81.260 26.370 81.790 ;
        RECT 25.355 81.230 26.355 81.260 ;
        RECT 25.355 81.000 26.355 81.020 ;
        RECT 22.000 80.700 23.150 80.790 ;
        RECT 25.330 80.700 26.370 81.000 ;
        RECT 26.530 80.960 26.850 81.290 ;
        RECT 22.000 80.560 26.370 80.700 ;
        RECT 22.000 80.540 25.380 80.560 ;
        RECT 18.690 79.620 23.010 79.890 ;
        RECT 15.345 79.130 16.345 79.160 ;
        RECT 15.345 78.900 16.345 78.920 ;
        RECT 15.330 78.600 16.370 78.900 ;
        RECT 16.520 78.860 18.550 79.190 ;
        RECT 18.690 79.070 19.690 79.620 ;
        RECT 19.870 79.160 20.130 79.190 ;
        RECT 18.690 78.900 19.690 78.910 ;
        RECT 18.690 78.690 19.700 78.900 ;
        RECT 19.850 78.870 20.130 79.160 ;
        RECT 19.870 78.850 20.130 78.870 ;
        RECT 18.550 78.600 19.700 78.690 ;
        RECT 15.330 78.460 19.700 78.600 ;
        RECT 16.320 78.440 19.700 78.460 ;
        RECT 14.250 77.590 16.370 77.860 ;
        RECT 14.250 75.760 14.600 77.590 ;
        RECT 14.850 76.760 15.170 77.090 ;
        RECT 15.330 77.060 16.360 77.590 ;
        RECT 17.090 77.090 17.820 78.440 ;
        RECT 20.380 77.790 21.320 79.620 ;
        RECT 21.570 79.160 21.830 79.190 ;
        RECT 21.570 78.870 21.850 79.160 ;
        RECT 22.010 79.070 23.010 79.620 ;
        RECT 23.880 79.190 24.610 80.540 ;
        RECT 27.100 79.960 27.450 81.790 ;
        RECT 25.330 79.690 27.450 79.960 ;
        RECT 22.010 78.900 23.010 78.910 ;
        RECT 21.570 78.850 21.830 78.870 ;
        RECT 22.000 78.690 23.010 78.900 ;
        RECT 23.150 78.860 25.180 79.190 ;
        RECT 25.340 79.160 26.370 79.690 ;
        RECT 25.355 79.130 26.355 79.160 ;
        RECT 25.355 78.900 26.355 78.920 ;
        RECT 22.000 78.600 23.150 78.690 ;
        RECT 25.330 78.600 26.370 78.900 ;
        RECT 26.530 78.860 26.850 79.190 ;
        RECT 22.000 78.460 26.370 78.600 ;
        RECT 22.000 78.440 25.380 78.460 ;
        RECT 18.690 77.520 23.010 77.790 ;
        RECT 15.345 77.030 16.345 77.060 ;
        RECT 15.345 76.800 16.345 76.820 ;
        RECT 15.330 76.500 16.370 76.800 ;
        RECT 16.520 76.760 18.550 77.090 ;
        RECT 18.690 76.970 19.690 77.520 ;
        RECT 19.870 77.060 20.130 77.090 ;
        RECT 18.690 76.800 19.690 76.810 ;
        RECT 18.690 76.590 19.700 76.800 ;
        RECT 19.850 76.770 20.130 77.060 ;
        RECT 19.870 76.750 20.130 76.770 ;
        RECT 18.550 76.500 19.700 76.590 ;
        RECT 15.330 76.360 19.700 76.500 ;
        RECT 16.320 76.340 19.700 76.360 ;
        RECT 14.250 75.490 16.370 75.760 ;
        RECT 14.250 73.660 14.600 75.490 ;
        RECT 14.850 74.660 15.170 74.990 ;
        RECT 15.330 74.960 16.360 75.490 ;
        RECT 17.090 74.990 17.820 76.340 ;
        RECT 20.380 75.690 21.320 77.520 ;
        RECT 21.570 77.060 21.830 77.090 ;
        RECT 21.570 76.770 21.850 77.060 ;
        RECT 22.010 76.970 23.010 77.520 ;
        RECT 23.880 77.090 24.610 78.440 ;
        RECT 27.100 77.860 27.450 79.690 ;
        RECT 25.330 77.590 27.450 77.860 ;
        RECT 22.010 76.800 23.010 76.810 ;
        RECT 21.570 76.750 21.830 76.770 ;
        RECT 22.000 76.590 23.010 76.800 ;
        RECT 23.150 76.760 25.180 77.090 ;
        RECT 25.340 77.060 26.370 77.590 ;
        RECT 25.355 77.030 26.355 77.060 ;
        RECT 25.355 76.800 26.355 76.820 ;
        RECT 22.000 76.500 23.150 76.590 ;
        RECT 25.330 76.500 26.370 76.800 ;
        RECT 26.530 76.760 26.850 77.090 ;
        RECT 22.000 76.360 26.370 76.500 ;
        RECT 22.000 76.340 25.380 76.360 ;
        RECT 18.690 75.420 23.010 75.690 ;
        RECT 15.345 74.930 16.345 74.960 ;
        RECT 15.345 74.700 16.345 74.720 ;
        RECT 15.330 74.400 16.370 74.700 ;
        RECT 16.520 74.660 18.550 74.990 ;
        RECT 18.690 74.870 19.690 75.420 ;
        RECT 19.870 74.960 20.130 74.990 ;
        RECT 18.690 74.700 19.690 74.710 ;
        RECT 18.690 74.490 19.700 74.700 ;
        RECT 19.850 74.670 20.130 74.960 ;
        RECT 19.870 74.650 20.130 74.670 ;
        RECT 18.550 74.400 19.700 74.490 ;
        RECT 15.330 74.260 19.700 74.400 ;
        RECT 16.320 74.240 19.700 74.260 ;
        RECT 14.250 73.390 16.370 73.660 ;
        RECT 14.250 71.560 14.600 73.390 ;
        RECT 14.850 72.560 15.170 72.890 ;
        RECT 15.330 72.860 16.360 73.390 ;
        RECT 17.090 72.890 17.820 74.240 ;
        RECT 20.380 73.590 21.320 75.420 ;
        RECT 21.570 74.960 21.830 74.990 ;
        RECT 21.570 74.670 21.850 74.960 ;
        RECT 22.010 74.870 23.010 75.420 ;
        RECT 23.880 74.990 24.610 76.340 ;
        RECT 27.100 75.760 27.450 77.590 ;
        RECT 25.330 75.490 27.450 75.760 ;
        RECT 22.010 74.700 23.010 74.710 ;
        RECT 21.570 74.650 21.830 74.670 ;
        RECT 22.000 74.490 23.010 74.700 ;
        RECT 23.150 74.660 25.180 74.990 ;
        RECT 25.340 74.960 26.370 75.490 ;
        RECT 25.355 74.930 26.355 74.960 ;
        RECT 25.355 74.700 26.355 74.720 ;
        RECT 22.000 74.400 23.150 74.490 ;
        RECT 25.330 74.400 26.370 74.700 ;
        RECT 26.530 74.660 26.850 74.990 ;
        RECT 22.000 74.260 26.370 74.400 ;
        RECT 22.000 74.240 25.380 74.260 ;
        RECT 18.690 73.320 23.010 73.590 ;
        RECT 15.345 72.830 16.345 72.860 ;
        RECT 15.345 72.600 16.345 72.620 ;
        RECT 15.330 72.300 16.370 72.600 ;
        RECT 16.520 72.560 18.550 72.890 ;
        RECT 18.690 72.770 19.690 73.320 ;
        RECT 19.870 72.860 20.130 72.890 ;
        RECT 18.690 72.600 19.690 72.610 ;
        RECT 18.690 72.390 19.700 72.600 ;
        RECT 19.850 72.570 20.130 72.860 ;
        RECT 19.870 72.550 20.130 72.570 ;
        RECT 18.550 72.300 19.700 72.390 ;
        RECT 15.330 72.160 19.700 72.300 ;
        RECT 16.320 72.140 19.700 72.160 ;
        RECT 14.250 71.290 16.370 71.560 ;
        RECT 14.250 69.460 14.600 71.290 ;
        RECT 14.850 70.460 15.170 70.790 ;
        RECT 15.330 70.760 16.360 71.290 ;
        RECT 17.090 70.790 17.820 72.140 ;
        RECT 20.380 71.490 21.320 73.320 ;
        RECT 21.570 72.860 21.830 72.890 ;
        RECT 21.570 72.570 21.850 72.860 ;
        RECT 22.010 72.770 23.010 73.320 ;
        RECT 23.880 72.890 24.610 74.240 ;
        RECT 27.100 73.660 27.450 75.490 ;
        RECT 25.330 73.390 27.450 73.660 ;
        RECT 22.010 72.600 23.010 72.610 ;
        RECT 21.570 72.550 21.830 72.570 ;
        RECT 22.000 72.390 23.010 72.600 ;
        RECT 23.150 72.560 25.180 72.890 ;
        RECT 25.340 72.860 26.370 73.390 ;
        RECT 25.355 72.830 26.355 72.860 ;
        RECT 25.355 72.600 26.355 72.620 ;
        RECT 22.000 72.300 23.150 72.390 ;
        RECT 25.330 72.300 26.370 72.600 ;
        RECT 26.530 72.560 26.850 72.890 ;
        RECT 22.000 72.160 26.370 72.300 ;
        RECT 22.000 72.140 25.380 72.160 ;
        RECT 18.690 71.220 23.010 71.490 ;
        RECT 15.345 70.730 16.345 70.760 ;
        RECT 15.345 70.500 16.345 70.520 ;
        RECT 15.330 70.200 16.370 70.500 ;
        RECT 16.520 70.460 18.550 70.790 ;
        RECT 18.690 70.670 19.690 71.220 ;
        RECT 19.870 70.760 20.130 70.790 ;
        RECT 18.690 70.500 19.690 70.510 ;
        RECT 18.690 70.290 19.700 70.500 ;
        RECT 19.850 70.470 20.130 70.760 ;
        RECT 19.870 70.450 20.130 70.470 ;
        RECT 18.550 70.200 19.700 70.290 ;
        RECT 15.330 70.060 19.700 70.200 ;
        RECT 16.320 70.040 19.700 70.060 ;
        RECT 14.250 69.190 16.370 69.460 ;
        RECT 14.250 67.360 14.600 69.190 ;
        RECT 14.850 68.360 15.170 68.690 ;
        RECT 15.330 68.660 16.360 69.190 ;
        RECT 17.090 68.690 17.820 70.040 ;
        RECT 20.380 69.390 21.320 71.220 ;
        RECT 21.570 70.760 21.830 70.790 ;
        RECT 21.570 70.470 21.850 70.760 ;
        RECT 22.010 70.670 23.010 71.220 ;
        RECT 23.880 70.790 24.610 72.140 ;
        RECT 27.100 71.560 27.450 73.390 ;
        RECT 25.330 71.290 27.450 71.560 ;
        RECT 22.010 70.500 23.010 70.510 ;
        RECT 21.570 70.450 21.830 70.470 ;
        RECT 22.000 70.290 23.010 70.500 ;
        RECT 23.150 70.460 25.180 70.790 ;
        RECT 25.340 70.760 26.370 71.290 ;
        RECT 25.355 70.730 26.355 70.760 ;
        RECT 25.355 70.500 26.355 70.520 ;
        RECT 22.000 70.200 23.150 70.290 ;
        RECT 25.330 70.200 26.370 70.500 ;
        RECT 26.530 70.460 26.850 70.790 ;
        RECT 22.000 70.060 26.370 70.200 ;
        RECT 22.000 70.040 25.380 70.060 ;
        RECT 18.690 69.120 23.010 69.390 ;
        RECT 15.345 68.630 16.345 68.660 ;
        RECT 15.345 68.400 16.345 68.420 ;
        RECT 15.330 68.100 16.370 68.400 ;
        RECT 16.520 68.360 18.550 68.690 ;
        RECT 18.690 68.570 19.690 69.120 ;
        RECT 19.870 68.660 20.130 68.690 ;
        RECT 18.690 68.400 19.690 68.410 ;
        RECT 18.690 68.190 19.700 68.400 ;
        RECT 19.850 68.370 20.130 68.660 ;
        RECT 19.870 68.350 20.130 68.370 ;
        RECT 18.550 68.100 19.700 68.190 ;
        RECT 15.330 67.960 19.700 68.100 ;
        RECT 16.320 67.940 19.700 67.960 ;
        RECT 14.250 67.090 16.370 67.360 ;
        RECT 14.250 65.260 14.600 67.090 ;
        RECT 14.850 66.260 15.170 66.590 ;
        RECT 15.330 66.560 16.360 67.090 ;
        RECT 17.090 66.590 17.820 67.940 ;
        RECT 20.380 67.290 21.320 69.120 ;
        RECT 21.570 68.660 21.830 68.690 ;
        RECT 21.570 68.370 21.850 68.660 ;
        RECT 22.010 68.570 23.010 69.120 ;
        RECT 23.880 68.690 24.610 70.040 ;
        RECT 27.100 69.460 27.450 71.290 ;
        RECT 25.330 69.190 27.450 69.460 ;
        RECT 22.010 68.400 23.010 68.410 ;
        RECT 21.570 68.350 21.830 68.370 ;
        RECT 22.000 68.190 23.010 68.400 ;
        RECT 23.150 68.360 25.180 68.690 ;
        RECT 25.340 68.660 26.370 69.190 ;
        RECT 25.355 68.630 26.355 68.660 ;
        RECT 25.355 68.400 26.355 68.420 ;
        RECT 22.000 68.100 23.150 68.190 ;
        RECT 25.330 68.100 26.370 68.400 ;
        RECT 26.530 68.360 26.850 68.690 ;
        RECT 22.000 67.960 26.370 68.100 ;
        RECT 22.000 67.940 25.380 67.960 ;
        RECT 18.690 67.020 23.010 67.290 ;
        RECT 15.345 66.530 16.345 66.560 ;
        RECT 15.345 66.300 16.345 66.320 ;
        RECT 15.330 66.000 16.370 66.300 ;
        RECT 16.520 66.260 18.550 66.590 ;
        RECT 18.690 66.470 19.690 67.020 ;
        RECT 19.870 66.560 20.130 66.590 ;
        RECT 18.690 66.300 19.690 66.310 ;
        RECT 18.690 66.090 19.700 66.300 ;
        RECT 19.850 66.270 20.130 66.560 ;
        RECT 19.870 66.250 20.130 66.270 ;
        RECT 18.550 66.000 19.700 66.090 ;
        RECT 15.330 65.860 19.700 66.000 ;
        RECT 16.320 65.840 19.700 65.860 ;
        RECT 14.250 64.990 16.370 65.260 ;
        RECT 14.250 63.160 14.600 64.990 ;
        RECT 14.850 64.160 15.170 64.490 ;
        RECT 15.330 64.460 16.360 64.990 ;
        RECT 17.090 64.490 17.820 65.840 ;
        RECT 20.380 65.190 21.320 67.020 ;
        RECT 21.570 66.560 21.830 66.590 ;
        RECT 21.570 66.270 21.850 66.560 ;
        RECT 22.010 66.470 23.010 67.020 ;
        RECT 23.880 66.590 24.610 67.940 ;
        RECT 27.100 67.360 27.450 69.190 ;
        RECT 25.330 67.090 27.450 67.360 ;
        RECT 22.010 66.300 23.010 66.310 ;
        RECT 21.570 66.250 21.830 66.270 ;
        RECT 22.000 66.090 23.010 66.300 ;
        RECT 23.150 66.260 25.180 66.590 ;
        RECT 25.340 66.560 26.370 67.090 ;
        RECT 25.355 66.530 26.355 66.560 ;
        RECT 25.355 66.300 26.355 66.320 ;
        RECT 22.000 66.000 23.150 66.090 ;
        RECT 25.330 66.000 26.370 66.300 ;
        RECT 26.530 66.260 26.850 66.590 ;
        RECT 22.000 65.860 26.370 66.000 ;
        RECT 22.000 65.840 25.380 65.860 ;
        RECT 18.690 64.920 23.010 65.190 ;
        RECT 15.345 64.430 16.345 64.460 ;
        RECT 15.345 64.200 16.345 64.220 ;
        RECT 15.330 63.900 16.370 64.200 ;
        RECT 16.520 64.160 18.550 64.490 ;
        RECT 18.690 64.370 19.690 64.920 ;
        RECT 19.870 64.460 20.130 64.490 ;
        RECT 18.690 64.200 19.690 64.210 ;
        RECT 18.690 63.990 19.700 64.200 ;
        RECT 19.850 64.170 20.130 64.460 ;
        RECT 19.870 64.150 20.130 64.170 ;
        RECT 18.550 63.900 19.700 63.990 ;
        RECT 15.330 63.760 19.700 63.900 ;
        RECT 16.320 63.740 19.700 63.760 ;
        RECT 14.250 62.890 16.370 63.160 ;
        RECT 14.250 61.060 14.600 62.890 ;
        RECT 14.850 62.060 15.170 62.390 ;
        RECT 15.330 62.360 16.360 62.890 ;
        RECT 17.090 62.390 17.820 63.740 ;
        RECT 20.380 63.090 21.320 64.920 ;
        RECT 21.570 64.460 21.830 64.490 ;
        RECT 21.570 64.170 21.850 64.460 ;
        RECT 22.010 64.370 23.010 64.920 ;
        RECT 23.880 64.490 24.610 65.840 ;
        RECT 27.100 65.260 27.450 67.090 ;
        RECT 25.330 64.990 27.450 65.260 ;
        RECT 22.010 64.200 23.010 64.210 ;
        RECT 21.570 64.150 21.830 64.170 ;
        RECT 22.000 63.990 23.010 64.200 ;
        RECT 23.150 64.160 25.180 64.490 ;
        RECT 25.340 64.460 26.370 64.990 ;
        RECT 25.355 64.430 26.355 64.460 ;
        RECT 25.355 64.200 26.355 64.220 ;
        RECT 22.000 63.900 23.150 63.990 ;
        RECT 25.330 63.900 26.370 64.200 ;
        RECT 26.530 64.160 26.850 64.490 ;
        RECT 22.000 63.760 26.370 63.900 ;
        RECT 22.000 63.740 25.380 63.760 ;
        RECT 18.690 62.820 23.010 63.090 ;
        RECT 15.345 62.330 16.345 62.360 ;
        RECT 15.345 62.100 16.345 62.120 ;
        RECT 15.330 61.800 16.370 62.100 ;
        RECT 16.520 62.060 18.550 62.390 ;
        RECT 18.690 62.270 19.690 62.820 ;
        RECT 19.870 62.360 20.130 62.390 ;
        RECT 18.690 62.100 19.690 62.110 ;
        RECT 18.690 61.890 19.700 62.100 ;
        RECT 19.850 62.070 20.130 62.360 ;
        RECT 19.870 62.050 20.130 62.070 ;
        RECT 18.550 61.800 19.700 61.890 ;
        RECT 15.330 61.660 19.700 61.800 ;
        RECT 16.320 61.640 19.700 61.660 ;
        RECT 14.250 60.790 16.370 61.060 ;
        RECT 14.250 58.960 14.600 60.790 ;
        RECT 14.850 59.960 15.170 60.290 ;
        RECT 15.330 60.260 16.360 60.790 ;
        RECT 17.090 60.290 17.820 61.640 ;
        RECT 20.380 60.990 21.320 62.820 ;
        RECT 21.570 62.360 21.830 62.390 ;
        RECT 21.570 62.070 21.850 62.360 ;
        RECT 22.010 62.270 23.010 62.820 ;
        RECT 23.880 62.390 24.610 63.740 ;
        RECT 27.100 63.160 27.450 64.990 ;
        RECT 25.330 62.890 27.450 63.160 ;
        RECT 22.010 62.100 23.010 62.110 ;
        RECT 21.570 62.050 21.830 62.070 ;
        RECT 22.000 61.890 23.010 62.100 ;
        RECT 23.150 62.060 25.180 62.390 ;
        RECT 25.340 62.360 26.370 62.890 ;
        RECT 25.355 62.330 26.355 62.360 ;
        RECT 25.355 62.100 26.355 62.120 ;
        RECT 22.000 61.800 23.150 61.890 ;
        RECT 25.330 61.800 26.370 62.100 ;
        RECT 26.530 62.060 26.850 62.390 ;
        RECT 22.000 61.660 26.370 61.800 ;
        RECT 22.000 61.640 25.380 61.660 ;
        RECT 18.690 60.720 23.010 60.990 ;
        RECT 15.345 60.230 16.345 60.260 ;
        RECT 15.345 60.000 16.345 60.020 ;
        RECT 15.330 59.700 16.370 60.000 ;
        RECT 16.520 59.960 18.550 60.290 ;
        RECT 18.690 60.170 19.690 60.720 ;
        RECT 19.870 60.260 20.130 60.290 ;
        RECT 18.690 60.000 19.690 60.010 ;
        RECT 18.690 59.790 19.700 60.000 ;
        RECT 19.850 59.970 20.130 60.260 ;
        RECT 19.870 59.950 20.130 59.970 ;
        RECT 18.550 59.700 19.700 59.790 ;
        RECT 15.330 59.560 19.700 59.700 ;
        RECT 16.320 59.540 19.700 59.560 ;
        RECT 14.250 58.690 16.370 58.960 ;
        RECT 14.250 56.860 14.600 58.690 ;
        RECT 14.850 57.860 15.170 58.190 ;
        RECT 15.330 58.160 16.360 58.690 ;
        RECT 17.090 58.190 17.820 59.540 ;
        RECT 20.380 58.890 21.320 60.720 ;
        RECT 21.570 60.260 21.830 60.290 ;
        RECT 21.570 59.970 21.850 60.260 ;
        RECT 22.010 60.170 23.010 60.720 ;
        RECT 23.880 60.290 24.610 61.640 ;
        RECT 27.100 61.060 27.450 62.890 ;
        RECT 25.330 60.790 27.450 61.060 ;
        RECT 22.010 60.000 23.010 60.010 ;
        RECT 21.570 59.950 21.830 59.970 ;
        RECT 22.000 59.790 23.010 60.000 ;
        RECT 23.150 59.960 25.180 60.290 ;
        RECT 25.340 60.260 26.370 60.790 ;
        RECT 25.355 60.230 26.355 60.260 ;
        RECT 25.355 60.000 26.355 60.020 ;
        RECT 22.000 59.700 23.150 59.790 ;
        RECT 25.330 59.700 26.370 60.000 ;
        RECT 26.530 59.960 26.850 60.290 ;
        RECT 22.000 59.560 26.370 59.700 ;
        RECT 22.000 59.540 25.380 59.560 ;
        RECT 18.690 58.620 23.010 58.890 ;
        RECT 15.345 58.130 16.345 58.160 ;
        RECT 15.345 57.900 16.345 57.920 ;
        RECT 15.330 57.600 16.370 57.900 ;
        RECT 16.520 57.860 18.550 58.190 ;
        RECT 18.690 58.070 19.690 58.620 ;
        RECT 19.870 58.160 20.130 58.190 ;
        RECT 18.690 57.900 19.690 57.910 ;
        RECT 18.690 57.690 19.700 57.900 ;
        RECT 19.850 57.870 20.130 58.160 ;
        RECT 19.870 57.850 20.130 57.870 ;
        RECT 18.550 57.600 19.700 57.690 ;
        RECT 15.330 57.460 19.700 57.600 ;
        RECT 16.320 57.440 19.700 57.460 ;
        RECT 14.250 56.590 16.370 56.860 ;
        RECT 14.250 54.760 14.600 56.590 ;
        RECT 14.850 55.760 15.170 56.090 ;
        RECT 15.330 56.060 16.360 56.590 ;
        RECT 17.090 56.090 17.820 57.440 ;
        RECT 20.380 56.790 21.320 58.620 ;
        RECT 21.570 58.160 21.830 58.190 ;
        RECT 21.570 57.870 21.850 58.160 ;
        RECT 22.010 58.070 23.010 58.620 ;
        RECT 23.880 58.190 24.610 59.540 ;
        RECT 27.100 58.960 27.450 60.790 ;
        RECT 25.330 58.690 27.450 58.960 ;
        RECT 22.010 57.900 23.010 57.910 ;
        RECT 21.570 57.850 21.830 57.870 ;
        RECT 22.000 57.690 23.010 57.900 ;
        RECT 23.150 57.860 25.180 58.190 ;
        RECT 25.340 58.160 26.370 58.690 ;
        RECT 25.355 58.130 26.355 58.160 ;
        RECT 25.355 57.900 26.355 57.920 ;
        RECT 22.000 57.600 23.150 57.690 ;
        RECT 25.330 57.600 26.370 57.900 ;
        RECT 26.530 57.860 26.850 58.190 ;
        RECT 22.000 57.460 26.370 57.600 ;
        RECT 22.000 57.440 25.380 57.460 ;
        RECT 18.690 56.520 23.010 56.790 ;
        RECT 15.345 56.030 16.345 56.060 ;
        RECT 15.345 55.800 16.345 55.820 ;
        RECT 15.330 55.500 16.370 55.800 ;
        RECT 16.520 55.760 18.550 56.090 ;
        RECT 18.690 55.970 19.690 56.520 ;
        RECT 19.870 56.060 20.130 56.090 ;
        RECT 18.690 55.800 19.690 55.810 ;
        RECT 18.690 55.590 19.700 55.800 ;
        RECT 19.850 55.770 20.130 56.060 ;
        RECT 19.870 55.750 20.130 55.770 ;
        RECT 18.550 55.500 19.700 55.590 ;
        RECT 15.330 55.360 19.700 55.500 ;
        RECT 16.320 55.340 19.700 55.360 ;
        RECT 14.250 54.490 16.370 54.760 ;
        RECT 14.250 52.660 14.600 54.490 ;
        RECT 14.850 53.660 15.170 53.990 ;
        RECT 15.330 53.960 16.360 54.490 ;
        RECT 17.090 53.990 17.820 55.340 ;
        RECT 20.380 54.690 21.320 56.520 ;
        RECT 21.570 56.060 21.830 56.090 ;
        RECT 21.570 55.770 21.850 56.060 ;
        RECT 22.010 55.970 23.010 56.520 ;
        RECT 23.880 56.090 24.610 57.440 ;
        RECT 27.100 56.860 27.450 58.690 ;
        RECT 25.330 56.590 27.450 56.860 ;
        RECT 22.010 55.800 23.010 55.810 ;
        RECT 21.570 55.750 21.830 55.770 ;
        RECT 22.000 55.590 23.010 55.800 ;
        RECT 23.150 55.760 25.180 56.090 ;
        RECT 25.340 56.060 26.370 56.590 ;
        RECT 25.355 56.030 26.355 56.060 ;
        RECT 25.355 55.800 26.355 55.820 ;
        RECT 22.000 55.500 23.150 55.590 ;
        RECT 25.330 55.500 26.370 55.800 ;
        RECT 26.530 55.760 26.850 56.090 ;
        RECT 22.000 55.360 26.370 55.500 ;
        RECT 22.000 55.340 25.380 55.360 ;
        RECT 18.690 54.420 23.010 54.690 ;
        RECT 15.345 53.930 16.345 53.960 ;
        RECT 15.345 53.700 16.345 53.720 ;
        RECT 15.330 53.400 16.370 53.700 ;
        RECT 16.520 53.660 18.550 53.990 ;
        RECT 18.690 53.870 19.690 54.420 ;
        RECT 19.870 53.960 20.130 53.990 ;
        RECT 18.690 53.700 19.690 53.710 ;
        RECT 18.690 53.490 19.700 53.700 ;
        RECT 19.850 53.670 20.130 53.960 ;
        RECT 19.870 53.650 20.130 53.670 ;
        RECT 18.550 53.400 19.700 53.490 ;
        RECT 15.330 53.260 19.700 53.400 ;
        RECT 16.320 53.240 19.700 53.260 ;
        RECT 14.250 52.390 16.370 52.660 ;
        RECT 14.250 50.560 14.600 52.390 ;
        RECT 14.850 51.560 15.170 51.890 ;
        RECT 15.330 51.860 16.360 52.390 ;
        RECT 17.090 51.890 17.820 53.240 ;
        RECT 20.380 52.590 21.320 54.420 ;
        RECT 21.570 53.960 21.830 53.990 ;
        RECT 21.570 53.670 21.850 53.960 ;
        RECT 22.010 53.870 23.010 54.420 ;
        RECT 23.880 53.990 24.610 55.340 ;
        RECT 27.100 54.760 27.450 56.590 ;
        RECT 25.330 54.490 27.450 54.760 ;
        RECT 22.010 53.700 23.010 53.710 ;
        RECT 21.570 53.650 21.830 53.670 ;
        RECT 22.000 53.490 23.010 53.700 ;
        RECT 23.150 53.660 25.180 53.990 ;
        RECT 25.340 53.960 26.370 54.490 ;
        RECT 25.355 53.930 26.355 53.960 ;
        RECT 25.355 53.700 26.355 53.720 ;
        RECT 22.000 53.400 23.150 53.490 ;
        RECT 25.330 53.400 26.370 53.700 ;
        RECT 26.530 53.660 26.850 53.990 ;
        RECT 22.000 53.260 26.370 53.400 ;
        RECT 22.000 53.240 25.380 53.260 ;
        RECT 18.690 52.320 23.010 52.590 ;
        RECT 15.345 51.830 16.345 51.860 ;
        RECT 15.345 51.600 16.345 51.620 ;
        RECT 15.330 51.300 16.370 51.600 ;
        RECT 16.520 51.560 18.550 51.890 ;
        RECT 18.690 51.770 19.690 52.320 ;
        RECT 19.870 51.860 20.130 51.890 ;
        RECT 18.690 51.600 19.690 51.610 ;
        RECT 18.690 51.390 19.700 51.600 ;
        RECT 19.850 51.570 20.130 51.860 ;
        RECT 19.870 51.550 20.130 51.570 ;
        RECT 18.550 51.300 19.700 51.390 ;
        RECT 15.330 51.160 19.700 51.300 ;
        RECT 16.320 51.140 19.700 51.160 ;
        RECT 14.250 50.290 16.370 50.560 ;
        RECT 14.250 48.460 14.600 50.290 ;
        RECT 14.850 49.460 15.170 49.790 ;
        RECT 15.330 49.760 16.360 50.290 ;
        RECT 17.090 49.790 17.820 51.140 ;
        RECT 20.380 50.490 21.320 52.320 ;
        RECT 21.570 51.860 21.830 51.890 ;
        RECT 21.570 51.570 21.850 51.860 ;
        RECT 22.010 51.770 23.010 52.320 ;
        RECT 23.880 51.890 24.610 53.240 ;
        RECT 27.100 52.660 27.450 54.490 ;
        RECT 25.330 52.390 27.450 52.660 ;
        RECT 22.010 51.600 23.010 51.610 ;
        RECT 21.570 51.550 21.830 51.570 ;
        RECT 22.000 51.390 23.010 51.600 ;
        RECT 23.150 51.560 25.180 51.890 ;
        RECT 25.340 51.860 26.370 52.390 ;
        RECT 25.355 51.830 26.355 51.860 ;
        RECT 25.355 51.600 26.355 51.620 ;
        RECT 22.000 51.300 23.150 51.390 ;
        RECT 25.330 51.300 26.370 51.600 ;
        RECT 26.530 51.560 26.850 51.890 ;
        RECT 22.000 51.160 26.370 51.300 ;
        RECT 22.000 51.140 25.380 51.160 ;
        RECT 18.690 50.220 23.010 50.490 ;
        RECT 15.345 49.730 16.345 49.760 ;
        RECT 15.345 49.500 16.345 49.520 ;
        RECT 15.330 49.200 16.370 49.500 ;
        RECT 16.520 49.460 18.550 49.790 ;
        RECT 18.690 49.670 19.690 50.220 ;
        RECT 19.870 49.760 20.130 49.790 ;
        RECT 18.690 49.500 19.690 49.510 ;
        RECT 18.690 49.290 19.700 49.500 ;
        RECT 19.850 49.470 20.130 49.760 ;
        RECT 19.870 49.450 20.130 49.470 ;
        RECT 18.550 49.200 19.700 49.290 ;
        RECT 15.330 49.060 19.700 49.200 ;
        RECT 16.320 49.040 19.700 49.060 ;
        RECT 14.250 48.190 16.370 48.460 ;
        RECT 14.250 46.360 14.600 48.190 ;
        RECT 14.850 47.360 15.170 47.690 ;
        RECT 15.330 47.660 16.360 48.190 ;
        RECT 17.090 47.690 17.820 49.040 ;
        RECT 20.380 48.390 21.320 50.220 ;
        RECT 21.570 49.760 21.830 49.790 ;
        RECT 21.570 49.470 21.850 49.760 ;
        RECT 22.010 49.670 23.010 50.220 ;
        RECT 23.880 49.790 24.610 51.140 ;
        RECT 27.100 50.560 27.450 52.390 ;
        RECT 25.330 50.290 27.450 50.560 ;
        RECT 22.010 49.500 23.010 49.510 ;
        RECT 21.570 49.450 21.830 49.470 ;
        RECT 22.000 49.290 23.010 49.500 ;
        RECT 23.150 49.460 25.180 49.790 ;
        RECT 25.340 49.760 26.370 50.290 ;
        RECT 25.355 49.730 26.355 49.760 ;
        RECT 25.355 49.500 26.355 49.520 ;
        RECT 22.000 49.200 23.150 49.290 ;
        RECT 25.330 49.200 26.370 49.500 ;
        RECT 26.530 49.460 26.850 49.790 ;
        RECT 22.000 49.060 26.370 49.200 ;
        RECT 22.000 49.040 25.380 49.060 ;
        RECT 18.690 48.120 23.010 48.390 ;
        RECT 15.345 47.630 16.345 47.660 ;
        RECT 15.345 47.400 16.345 47.420 ;
        RECT 15.330 47.100 16.370 47.400 ;
        RECT 16.520 47.360 18.550 47.690 ;
        RECT 18.690 47.570 19.690 48.120 ;
        RECT 19.870 47.660 20.130 47.690 ;
        RECT 18.690 47.400 19.690 47.410 ;
        RECT 18.690 47.190 19.700 47.400 ;
        RECT 19.850 47.370 20.130 47.660 ;
        RECT 19.870 47.350 20.130 47.370 ;
        RECT 18.550 47.100 19.700 47.190 ;
        RECT 15.330 46.960 19.700 47.100 ;
        RECT 16.320 46.940 19.700 46.960 ;
        RECT 14.250 46.090 16.370 46.360 ;
        RECT 14.250 44.260 14.600 46.090 ;
        RECT 14.850 45.260 15.170 45.590 ;
        RECT 15.330 45.560 16.360 46.090 ;
        RECT 17.090 45.590 17.820 46.940 ;
        RECT 20.380 46.290 21.320 48.120 ;
        RECT 21.570 47.660 21.830 47.690 ;
        RECT 21.570 47.370 21.850 47.660 ;
        RECT 22.010 47.570 23.010 48.120 ;
        RECT 23.880 47.690 24.610 49.040 ;
        RECT 27.100 48.460 27.450 50.290 ;
        RECT 25.330 48.190 27.450 48.460 ;
        RECT 22.010 47.400 23.010 47.410 ;
        RECT 21.570 47.350 21.830 47.370 ;
        RECT 22.000 47.190 23.010 47.400 ;
        RECT 23.150 47.360 25.180 47.690 ;
        RECT 25.340 47.660 26.370 48.190 ;
        RECT 25.355 47.630 26.355 47.660 ;
        RECT 25.355 47.400 26.355 47.420 ;
        RECT 22.000 47.100 23.150 47.190 ;
        RECT 25.330 47.100 26.370 47.400 ;
        RECT 26.530 47.360 26.850 47.690 ;
        RECT 22.000 46.960 26.370 47.100 ;
        RECT 22.000 46.940 25.380 46.960 ;
        RECT 18.690 46.020 23.010 46.290 ;
        RECT 15.345 45.530 16.345 45.560 ;
        RECT 15.345 45.300 16.345 45.320 ;
        RECT 15.330 45.000 16.370 45.300 ;
        RECT 16.520 45.260 18.550 45.590 ;
        RECT 18.690 45.470 19.690 46.020 ;
        RECT 19.870 45.560 20.130 45.590 ;
        RECT 18.690 45.300 19.690 45.310 ;
        RECT 18.690 45.090 19.700 45.300 ;
        RECT 19.850 45.270 20.130 45.560 ;
        RECT 19.870 45.250 20.130 45.270 ;
        RECT 18.550 45.000 19.700 45.090 ;
        RECT 15.330 44.860 19.700 45.000 ;
        RECT 16.320 44.840 19.700 44.860 ;
        RECT 14.250 43.990 16.370 44.260 ;
        RECT 14.250 42.160 14.600 43.990 ;
        RECT 14.850 43.160 15.170 43.490 ;
        RECT 15.330 43.460 16.360 43.990 ;
        RECT 17.090 43.490 17.820 44.840 ;
        RECT 20.380 44.190 21.320 46.020 ;
        RECT 21.570 45.560 21.830 45.590 ;
        RECT 21.570 45.270 21.850 45.560 ;
        RECT 22.010 45.470 23.010 46.020 ;
        RECT 23.880 45.590 24.610 46.940 ;
        RECT 27.100 46.360 27.450 48.190 ;
        RECT 25.330 46.090 27.450 46.360 ;
        RECT 22.010 45.300 23.010 45.310 ;
        RECT 21.570 45.250 21.830 45.270 ;
        RECT 22.000 45.090 23.010 45.300 ;
        RECT 23.150 45.260 25.180 45.590 ;
        RECT 25.340 45.560 26.370 46.090 ;
        RECT 25.355 45.530 26.355 45.560 ;
        RECT 25.355 45.300 26.355 45.320 ;
        RECT 22.000 45.000 23.150 45.090 ;
        RECT 25.330 45.000 26.370 45.300 ;
        RECT 26.530 45.260 26.850 45.590 ;
        RECT 22.000 44.860 26.370 45.000 ;
        RECT 22.000 44.840 25.380 44.860 ;
        RECT 18.690 43.920 23.010 44.190 ;
        RECT 15.345 43.430 16.345 43.460 ;
        RECT 15.345 43.200 16.345 43.220 ;
        RECT 15.330 42.900 16.370 43.200 ;
        RECT 16.520 43.160 18.550 43.490 ;
        RECT 18.690 43.370 19.690 43.920 ;
        RECT 19.870 43.460 20.130 43.490 ;
        RECT 18.690 43.200 19.690 43.210 ;
        RECT 18.690 42.990 19.700 43.200 ;
        RECT 19.850 43.170 20.130 43.460 ;
        RECT 19.870 43.150 20.130 43.170 ;
        RECT 18.550 42.900 19.700 42.990 ;
        RECT 15.330 42.760 19.700 42.900 ;
        RECT 16.320 42.740 19.700 42.760 ;
        RECT 14.250 41.890 16.370 42.160 ;
        RECT 14.250 40.060 14.600 41.890 ;
        RECT 14.850 41.060 15.170 41.390 ;
        RECT 15.330 41.360 16.360 41.890 ;
        RECT 17.090 41.390 17.820 42.740 ;
        RECT 20.380 42.090 21.320 43.920 ;
        RECT 21.570 43.460 21.830 43.490 ;
        RECT 21.570 43.170 21.850 43.460 ;
        RECT 22.010 43.370 23.010 43.920 ;
        RECT 23.880 43.490 24.610 44.840 ;
        RECT 27.100 44.260 27.450 46.090 ;
        RECT 25.330 43.990 27.450 44.260 ;
        RECT 22.010 43.200 23.010 43.210 ;
        RECT 21.570 43.150 21.830 43.170 ;
        RECT 22.000 42.990 23.010 43.200 ;
        RECT 23.150 43.160 25.180 43.490 ;
        RECT 25.340 43.460 26.370 43.990 ;
        RECT 25.355 43.430 26.355 43.460 ;
        RECT 25.355 43.200 26.355 43.220 ;
        RECT 22.000 42.900 23.150 42.990 ;
        RECT 25.330 42.900 26.370 43.200 ;
        RECT 26.530 43.160 26.850 43.490 ;
        RECT 22.000 42.760 26.370 42.900 ;
        RECT 22.000 42.740 25.380 42.760 ;
        RECT 18.690 41.820 23.010 42.090 ;
        RECT 15.345 41.330 16.345 41.360 ;
        RECT 15.345 41.100 16.345 41.120 ;
        RECT 15.330 40.800 16.370 41.100 ;
        RECT 16.520 41.060 18.550 41.390 ;
        RECT 18.690 41.270 19.690 41.820 ;
        RECT 19.870 41.360 20.130 41.390 ;
        RECT 18.690 41.100 19.690 41.110 ;
        RECT 18.690 40.890 19.700 41.100 ;
        RECT 19.850 41.070 20.130 41.360 ;
        RECT 19.870 41.050 20.130 41.070 ;
        RECT 18.550 40.800 19.700 40.890 ;
        RECT 15.330 40.660 19.700 40.800 ;
        RECT 16.320 40.640 19.700 40.660 ;
        RECT 14.250 39.790 16.370 40.060 ;
        RECT 14.250 37.960 14.600 39.790 ;
        RECT 14.850 38.960 15.170 39.290 ;
        RECT 15.330 39.260 16.360 39.790 ;
        RECT 17.090 39.290 17.820 40.640 ;
        RECT 20.380 39.990 21.320 41.820 ;
        RECT 21.570 41.360 21.830 41.390 ;
        RECT 21.570 41.070 21.850 41.360 ;
        RECT 22.010 41.270 23.010 41.820 ;
        RECT 23.880 41.390 24.610 42.740 ;
        RECT 27.100 42.160 27.450 43.990 ;
        RECT 25.330 41.890 27.450 42.160 ;
        RECT 22.010 41.100 23.010 41.110 ;
        RECT 21.570 41.050 21.830 41.070 ;
        RECT 22.000 40.890 23.010 41.100 ;
        RECT 23.150 41.060 25.180 41.390 ;
        RECT 25.340 41.360 26.370 41.890 ;
        RECT 25.355 41.330 26.355 41.360 ;
        RECT 25.355 41.100 26.355 41.120 ;
        RECT 22.000 40.800 23.150 40.890 ;
        RECT 25.330 40.800 26.370 41.100 ;
        RECT 26.530 41.060 26.850 41.390 ;
        RECT 22.000 40.660 26.370 40.800 ;
        RECT 22.000 40.640 25.380 40.660 ;
        RECT 18.690 39.720 23.010 39.990 ;
        RECT 15.345 39.230 16.345 39.260 ;
        RECT 15.345 39.000 16.345 39.020 ;
        RECT 15.330 38.700 16.370 39.000 ;
        RECT 16.520 38.960 18.550 39.290 ;
        RECT 18.690 39.170 19.690 39.720 ;
        RECT 19.870 39.260 20.130 39.290 ;
        RECT 18.690 39.000 19.690 39.010 ;
        RECT 18.690 38.790 19.700 39.000 ;
        RECT 19.850 38.970 20.130 39.260 ;
        RECT 19.870 38.950 20.130 38.970 ;
        RECT 18.550 38.700 19.700 38.790 ;
        RECT 15.330 38.560 19.700 38.700 ;
        RECT 16.320 38.540 19.700 38.560 ;
        RECT 14.250 37.690 16.370 37.960 ;
        RECT 14.250 35.860 14.600 37.690 ;
        RECT 14.850 36.860 15.170 37.190 ;
        RECT 15.330 37.160 16.360 37.690 ;
        RECT 17.090 37.190 17.820 38.540 ;
        RECT 20.380 37.890 21.320 39.720 ;
        RECT 21.570 39.260 21.830 39.290 ;
        RECT 21.570 38.970 21.850 39.260 ;
        RECT 22.010 39.170 23.010 39.720 ;
        RECT 23.880 39.290 24.610 40.640 ;
        RECT 27.100 40.060 27.450 41.890 ;
        RECT 25.330 39.790 27.450 40.060 ;
        RECT 22.010 39.000 23.010 39.010 ;
        RECT 21.570 38.950 21.830 38.970 ;
        RECT 22.000 38.790 23.010 39.000 ;
        RECT 23.150 38.960 25.180 39.290 ;
        RECT 25.340 39.260 26.370 39.790 ;
        RECT 25.355 39.230 26.355 39.260 ;
        RECT 25.355 39.000 26.355 39.020 ;
        RECT 22.000 38.700 23.150 38.790 ;
        RECT 25.330 38.700 26.370 39.000 ;
        RECT 26.530 38.960 26.850 39.290 ;
        RECT 22.000 38.560 26.370 38.700 ;
        RECT 22.000 38.540 25.380 38.560 ;
        RECT 18.690 37.620 23.010 37.890 ;
        RECT 15.345 37.130 16.345 37.160 ;
        RECT 15.345 36.900 16.345 36.920 ;
        RECT 15.330 36.600 16.370 36.900 ;
        RECT 16.520 36.860 18.550 37.190 ;
        RECT 18.690 37.070 19.690 37.620 ;
        RECT 19.870 37.160 20.130 37.190 ;
        RECT 18.690 36.900 19.690 36.910 ;
        RECT 18.690 36.690 19.700 36.900 ;
        RECT 19.850 36.870 20.130 37.160 ;
        RECT 19.870 36.850 20.130 36.870 ;
        RECT 18.550 36.600 19.700 36.690 ;
        RECT 15.330 36.460 19.700 36.600 ;
        RECT 16.320 36.440 19.700 36.460 ;
        RECT 14.250 35.590 16.370 35.860 ;
        RECT 14.250 33.760 14.600 35.590 ;
        RECT 14.850 34.760 15.170 35.090 ;
        RECT 15.330 35.060 16.360 35.590 ;
        RECT 17.090 35.090 17.820 36.440 ;
        RECT 20.380 35.790 21.320 37.620 ;
        RECT 21.570 37.160 21.830 37.190 ;
        RECT 21.570 36.870 21.850 37.160 ;
        RECT 22.010 37.070 23.010 37.620 ;
        RECT 23.880 37.190 24.610 38.540 ;
        RECT 27.100 37.960 27.450 39.790 ;
        RECT 25.330 37.690 27.450 37.960 ;
        RECT 22.010 36.900 23.010 36.910 ;
        RECT 21.570 36.850 21.830 36.870 ;
        RECT 22.000 36.690 23.010 36.900 ;
        RECT 23.150 36.860 25.180 37.190 ;
        RECT 25.340 37.160 26.370 37.690 ;
        RECT 25.355 37.130 26.355 37.160 ;
        RECT 25.355 36.900 26.355 36.920 ;
        RECT 22.000 36.600 23.150 36.690 ;
        RECT 25.330 36.600 26.370 36.900 ;
        RECT 26.530 36.860 26.850 37.190 ;
        RECT 22.000 36.460 26.370 36.600 ;
        RECT 22.000 36.440 25.380 36.460 ;
        RECT 18.690 35.520 23.010 35.790 ;
        RECT 15.345 35.030 16.345 35.060 ;
        RECT 15.345 34.800 16.345 34.820 ;
        RECT 15.330 34.500 16.370 34.800 ;
        RECT 16.520 34.760 18.550 35.090 ;
        RECT 18.690 34.970 19.690 35.520 ;
        RECT 19.870 35.060 20.130 35.090 ;
        RECT 18.690 34.800 19.690 34.810 ;
        RECT 18.690 34.590 19.700 34.800 ;
        RECT 19.850 34.770 20.130 35.060 ;
        RECT 19.870 34.750 20.130 34.770 ;
        RECT 18.550 34.500 19.700 34.590 ;
        RECT 15.330 34.360 19.700 34.500 ;
        RECT 16.320 34.340 19.700 34.360 ;
        RECT 14.250 33.490 16.370 33.760 ;
        RECT 14.250 31.660 14.600 33.490 ;
        RECT 14.850 32.660 15.170 32.990 ;
        RECT 15.330 32.960 16.360 33.490 ;
        RECT 17.090 32.990 17.820 34.340 ;
        RECT 20.380 33.690 21.320 35.520 ;
        RECT 21.570 35.060 21.830 35.090 ;
        RECT 21.570 34.770 21.850 35.060 ;
        RECT 22.010 34.970 23.010 35.520 ;
        RECT 23.880 35.090 24.610 36.440 ;
        RECT 27.100 35.860 27.450 37.690 ;
        RECT 25.330 35.590 27.450 35.860 ;
        RECT 22.010 34.800 23.010 34.810 ;
        RECT 21.570 34.750 21.830 34.770 ;
        RECT 22.000 34.590 23.010 34.800 ;
        RECT 23.150 34.760 25.180 35.090 ;
        RECT 25.340 35.060 26.370 35.590 ;
        RECT 25.355 35.030 26.355 35.060 ;
        RECT 25.355 34.800 26.355 34.820 ;
        RECT 22.000 34.500 23.150 34.590 ;
        RECT 25.330 34.500 26.370 34.800 ;
        RECT 26.530 34.760 26.850 35.090 ;
        RECT 22.000 34.360 26.370 34.500 ;
        RECT 22.000 34.340 25.380 34.360 ;
        RECT 18.690 33.420 23.010 33.690 ;
        RECT 15.345 32.930 16.345 32.960 ;
        RECT 15.345 32.700 16.345 32.720 ;
        RECT 15.330 32.400 16.370 32.700 ;
        RECT 16.520 32.660 18.550 32.990 ;
        RECT 18.690 32.870 19.690 33.420 ;
        RECT 19.870 32.960 20.130 32.990 ;
        RECT 18.690 32.700 19.690 32.710 ;
        RECT 18.690 32.490 19.700 32.700 ;
        RECT 19.850 32.670 20.130 32.960 ;
        RECT 19.870 32.650 20.130 32.670 ;
        RECT 18.550 32.400 19.700 32.490 ;
        RECT 15.330 32.260 19.700 32.400 ;
        RECT 16.320 32.240 19.700 32.260 ;
        RECT 14.250 31.390 16.370 31.660 ;
        RECT 14.250 29.560 14.600 31.390 ;
        RECT 14.850 30.560 15.170 30.890 ;
        RECT 15.330 30.860 16.360 31.390 ;
        RECT 17.090 30.890 17.820 32.240 ;
        RECT 20.380 31.590 21.320 33.420 ;
        RECT 21.570 32.960 21.830 32.990 ;
        RECT 21.570 32.670 21.850 32.960 ;
        RECT 22.010 32.870 23.010 33.420 ;
        RECT 23.880 32.990 24.610 34.340 ;
        RECT 27.100 33.760 27.450 35.590 ;
        RECT 25.330 33.490 27.450 33.760 ;
        RECT 22.010 32.700 23.010 32.710 ;
        RECT 21.570 32.650 21.830 32.670 ;
        RECT 22.000 32.490 23.010 32.700 ;
        RECT 23.150 32.660 25.180 32.990 ;
        RECT 25.340 32.960 26.370 33.490 ;
        RECT 25.355 32.930 26.355 32.960 ;
        RECT 25.355 32.700 26.355 32.720 ;
        RECT 22.000 32.400 23.150 32.490 ;
        RECT 25.330 32.400 26.370 32.700 ;
        RECT 26.530 32.660 26.850 32.990 ;
        RECT 22.000 32.260 26.370 32.400 ;
        RECT 22.000 32.240 25.380 32.260 ;
        RECT 18.690 31.320 23.010 31.590 ;
        RECT 15.345 30.830 16.345 30.860 ;
        RECT 15.345 30.600 16.345 30.620 ;
        RECT 15.330 30.300 16.370 30.600 ;
        RECT 16.520 30.560 18.550 30.890 ;
        RECT 18.690 30.770 19.690 31.320 ;
        RECT 19.870 30.860 20.130 30.890 ;
        RECT 18.690 30.600 19.690 30.610 ;
        RECT 18.690 30.390 19.700 30.600 ;
        RECT 19.850 30.570 20.130 30.860 ;
        RECT 19.870 30.550 20.130 30.570 ;
        RECT 18.550 30.300 19.700 30.390 ;
        RECT 15.330 30.160 19.700 30.300 ;
        RECT 16.320 30.140 19.700 30.160 ;
        RECT 14.250 29.290 16.370 29.560 ;
        RECT 14.250 27.460 14.600 29.290 ;
        RECT 14.850 28.460 15.170 28.790 ;
        RECT 15.330 28.760 16.360 29.290 ;
        RECT 17.090 28.790 17.820 30.140 ;
        RECT 20.380 29.490 21.320 31.320 ;
        RECT 21.570 30.860 21.830 30.890 ;
        RECT 21.570 30.570 21.850 30.860 ;
        RECT 22.010 30.770 23.010 31.320 ;
        RECT 23.880 30.890 24.610 32.240 ;
        RECT 27.100 31.660 27.450 33.490 ;
        RECT 25.330 31.390 27.450 31.660 ;
        RECT 22.010 30.600 23.010 30.610 ;
        RECT 21.570 30.550 21.830 30.570 ;
        RECT 22.000 30.390 23.010 30.600 ;
        RECT 23.150 30.560 25.180 30.890 ;
        RECT 25.340 30.860 26.370 31.390 ;
        RECT 25.355 30.830 26.355 30.860 ;
        RECT 25.355 30.600 26.355 30.620 ;
        RECT 22.000 30.300 23.150 30.390 ;
        RECT 25.330 30.300 26.370 30.600 ;
        RECT 26.530 30.560 26.850 30.890 ;
        RECT 22.000 30.160 26.370 30.300 ;
        RECT 22.000 30.140 25.380 30.160 ;
        RECT 18.690 29.220 23.010 29.490 ;
        RECT 15.345 28.730 16.345 28.760 ;
        RECT 15.345 28.500 16.345 28.520 ;
        RECT 15.330 28.200 16.370 28.500 ;
        RECT 16.520 28.460 18.550 28.790 ;
        RECT 18.690 28.670 19.690 29.220 ;
        RECT 19.870 28.760 20.130 28.790 ;
        RECT 18.690 28.500 19.690 28.510 ;
        RECT 18.690 28.290 19.700 28.500 ;
        RECT 19.850 28.470 20.130 28.760 ;
        RECT 19.870 28.450 20.130 28.470 ;
        RECT 18.550 28.200 19.700 28.290 ;
        RECT 15.330 28.060 19.700 28.200 ;
        RECT 16.320 28.040 19.700 28.060 ;
        RECT 14.250 27.190 16.370 27.460 ;
        RECT 14.250 25.360 14.600 27.190 ;
        RECT 14.850 26.360 15.170 26.690 ;
        RECT 15.330 26.660 16.360 27.190 ;
        RECT 17.090 26.690 17.820 28.040 ;
        RECT 20.380 27.390 21.320 29.220 ;
        RECT 21.570 28.760 21.830 28.790 ;
        RECT 21.570 28.470 21.850 28.760 ;
        RECT 22.010 28.670 23.010 29.220 ;
        RECT 23.880 28.790 24.610 30.140 ;
        RECT 27.100 29.560 27.450 31.390 ;
        RECT 25.330 29.290 27.450 29.560 ;
        RECT 22.010 28.500 23.010 28.510 ;
        RECT 21.570 28.450 21.830 28.470 ;
        RECT 22.000 28.290 23.010 28.500 ;
        RECT 23.150 28.460 25.180 28.790 ;
        RECT 25.340 28.760 26.370 29.290 ;
        RECT 25.355 28.730 26.355 28.760 ;
        RECT 25.355 28.500 26.355 28.520 ;
        RECT 22.000 28.200 23.150 28.290 ;
        RECT 25.330 28.200 26.370 28.500 ;
        RECT 26.530 28.460 26.850 28.790 ;
        RECT 22.000 28.060 26.370 28.200 ;
        RECT 22.000 28.040 25.380 28.060 ;
        RECT 18.690 27.120 23.010 27.390 ;
        RECT 15.345 26.630 16.345 26.660 ;
        RECT 15.345 26.400 16.345 26.420 ;
        RECT 15.330 26.100 16.370 26.400 ;
        RECT 16.520 26.360 18.550 26.690 ;
        RECT 18.690 26.570 19.690 27.120 ;
        RECT 19.870 26.660 20.130 26.690 ;
        RECT 18.690 26.400 19.690 26.410 ;
        RECT 18.690 26.190 19.700 26.400 ;
        RECT 19.850 26.370 20.130 26.660 ;
        RECT 19.870 26.350 20.130 26.370 ;
        RECT 18.550 26.100 19.700 26.190 ;
        RECT 15.330 25.960 19.700 26.100 ;
        RECT 16.320 25.940 19.700 25.960 ;
        RECT 14.250 25.090 16.370 25.360 ;
        RECT 14.250 23.260 14.600 25.090 ;
        RECT 14.850 24.260 15.170 24.590 ;
        RECT 15.330 24.560 16.360 25.090 ;
        RECT 17.090 24.590 17.820 25.940 ;
        RECT 20.380 25.290 21.320 27.120 ;
        RECT 21.570 26.660 21.830 26.690 ;
        RECT 21.570 26.370 21.850 26.660 ;
        RECT 22.010 26.570 23.010 27.120 ;
        RECT 23.880 26.690 24.610 28.040 ;
        RECT 27.100 27.460 27.450 29.290 ;
        RECT 25.330 27.190 27.450 27.460 ;
        RECT 22.010 26.400 23.010 26.410 ;
        RECT 21.570 26.350 21.830 26.370 ;
        RECT 22.000 26.190 23.010 26.400 ;
        RECT 23.150 26.360 25.180 26.690 ;
        RECT 25.340 26.660 26.370 27.190 ;
        RECT 25.355 26.630 26.355 26.660 ;
        RECT 25.355 26.400 26.355 26.420 ;
        RECT 22.000 26.100 23.150 26.190 ;
        RECT 25.330 26.100 26.370 26.400 ;
        RECT 26.530 26.360 26.850 26.690 ;
        RECT 22.000 25.960 26.370 26.100 ;
        RECT 22.000 25.940 25.380 25.960 ;
        RECT 18.690 25.020 23.010 25.290 ;
        RECT 15.345 24.530 16.345 24.560 ;
        RECT 15.345 24.300 16.345 24.320 ;
        RECT 15.330 24.000 16.370 24.300 ;
        RECT 16.520 24.260 18.550 24.590 ;
        RECT 18.690 24.470 19.690 25.020 ;
        RECT 19.870 24.560 20.130 24.590 ;
        RECT 18.690 24.300 19.690 24.310 ;
        RECT 18.690 24.090 19.700 24.300 ;
        RECT 19.850 24.270 20.130 24.560 ;
        RECT 19.870 24.250 20.130 24.270 ;
        RECT 18.550 24.000 19.700 24.090 ;
        RECT 15.330 23.860 19.700 24.000 ;
        RECT 16.320 23.840 19.700 23.860 ;
        RECT 14.250 22.990 16.370 23.260 ;
        RECT 14.250 21.160 14.600 22.990 ;
        RECT 14.850 22.160 15.170 22.490 ;
        RECT 15.330 22.460 16.360 22.990 ;
        RECT 17.090 22.490 17.820 23.840 ;
        RECT 20.380 23.190 21.320 25.020 ;
        RECT 21.570 24.560 21.830 24.590 ;
        RECT 21.570 24.270 21.850 24.560 ;
        RECT 22.010 24.470 23.010 25.020 ;
        RECT 23.880 24.590 24.610 25.940 ;
        RECT 27.100 25.360 27.450 27.190 ;
        RECT 25.330 25.090 27.450 25.360 ;
        RECT 22.010 24.300 23.010 24.310 ;
        RECT 21.570 24.250 21.830 24.270 ;
        RECT 22.000 24.090 23.010 24.300 ;
        RECT 23.150 24.260 25.180 24.590 ;
        RECT 25.340 24.560 26.370 25.090 ;
        RECT 25.355 24.530 26.355 24.560 ;
        RECT 25.355 24.300 26.355 24.320 ;
        RECT 22.000 24.000 23.150 24.090 ;
        RECT 25.330 24.000 26.370 24.300 ;
        RECT 26.530 24.260 26.850 24.590 ;
        RECT 22.000 23.860 26.370 24.000 ;
        RECT 22.000 23.840 25.380 23.860 ;
        RECT 18.690 22.920 23.010 23.190 ;
        RECT 15.345 22.430 16.345 22.460 ;
        RECT 15.345 22.200 16.345 22.220 ;
        RECT 15.330 21.900 16.370 22.200 ;
        RECT 16.520 22.160 18.550 22.490 ;
        RECT 18.690 22.370 19.690 22.920 ;
        RECT 19.870 22.460 20.130 22.490 ;
        RECT 18.690 22.200 19.690 22.210 ;
        RECT 18.690 21.990 19.700 22.200 ;
        RECT 19.850 22.170 20.130 22.460 ;
        RECT 19.870 22.150 20.130 22.170 ;
        RECT 18.550 21.900 19.700 21.990 ;
        RECT 15.330 21.760 19.700 21.900 ;
        RECT 16.320 21.740 19.700 21.760 ;
        RECT 14.250 20.890 16.370 21.160 ;
        RECT 14.250 19.060 14.600 20.890 ;
        RECT 14.850 20.060 15.170 20.390 ;
        RECT 15.330 20.360 16.360 20.890 ;
        RECT 17.090 20.390 17.820 21.740 ;
        RECT 20.380 21.090 21.320 22.920 ;
        RECT 21.570 22.460 21.830 22.490 ;
        RECT 21.570 22.170 21.850 22.460 ;
        RECT 22.010 22.370 23.010 22.920 ;
        RECT 23.880 22.490 24.610 23.840 ;
        RECT 27.100 23.260 27.450 25.090 ;
        RECT 25.330 22.990 27.450 23.260 ;
        RECT 22.010 22.200 23.010 22.210 ;
        RECT 21.570 22.150 21.830 22.170 ;
        RECT 22.000 21.990 23.010 22.200 ;
        RECT 23.150 22.160 25.180 22.490 ;
        RECT 25.340 22.460 26.370 22.990 ;
        RECT 25.355 22.430 26.355 22.460 ;
        RECT 25.355 22.200 26.355 22.220 ;
        RECT 22.000 21.900 23.150 21.990 ;
        RECT 25.330 21.900 26.370 22.200 ;
        RECT 26.530 22.160 26.850 22.490 ;
        RECT 22.000 21.760 26.370 21.900 ;
        RECT 22.000 21.740 25.380 21.760 ;
        RECT 18.690 20.820 23.010 21.090 ;
        RECT 15.345 20.330 16.345 20.360 ;
        RECT 15.345 20.100 16.345 20.120 ;
        RECT 15.330 19.800 16.370 20.100 ;
        RECT 16.520 20.060 18.550 20.390 ;
        RECT 18.690 20.270 19.690 20.820 ;
        RECT 19.870 20.360 20.130 20.390 ;
        RECT 18.690 20.100 19.690 20.110 ;
        RECT 18.690 19.890 19.700 20.100 ;
        RECT 19.850 20.070 20.130 20.360 ;
        RECT 19.870 20.050 20.130 20.070 ;
        RECT 18.550 19.800 19.700 19.890 ;
        RECT 15.330 19.660 19.700 19.800 ;
        RECT 16.320 19.640 19.700 19.660 ;
        RECT 14.250 18.790 16.370 19.060 ;
        RECT 14.250 16.960 14.600 18.790 ;
        RECT 14.850 17.960 15.170 18.290 ;
        RECT 15.330 18.260 16.360 18.790 ;
        RECT 17.090 18.290 17.820 19.640 ;
        RECT 20.380 18.990 21.320 20.820 ;
        RECT 21.570 20.360 21.830 20.390 ;
        RECT 21.570 20.070 21.850 20.360 ;
        RECT 22.010 20.270 23.010 20.820 ;
        RECT 23.880 20.390 24.610 21.740 ;
        RECT 27.100 21.160 27.450 22.990 ;
        RECT 25.330 20.890 27.450 21.160 ;
        RECT 22.010 20.100 23.010 20.110 ;
        RECT 21.570 20.050 21.830 20.070 ;
        RECT 22.000 19.890 23.010 20.100 ;
        RECT 23.150 20.060 25.180 20.390 ;
        RECT 25.340 20.360 26.370 20.890 ;
        RECT 25.355 20.330 26.355 20.360 ;
        RECT 25.355 20.100 26.355 20.120 ;
        RECT 22.000 19.800 23.150 19.890 ;
        RECT 25.330 19.800 26.370 20.100 ;
        RECT 26.530 20.060 26.850 20.390 ;
        RECT 22.000 19.660 26.370 19.800 ;
        RECT 22.000 19.640 25.380 19.660 ;
        RECT 18.690 18.720 23.010 18.990 ;
        RECT 15.345 18.230 16.345 18.260 ;
        RECT 15.345 18.000 16.345 18.020 ;
        RECT 15.330 17.700 16.370 18.000 ;
        RECT 16.520 17.960 18.550 18.290 ;
        RECT 18.690 18.170 19.690 18.720 ;
        RECT 19.870 18.260 20.130 18.290 ;
        RECT 18.690 18.000 19.690 18.010 ;
        RECT 18.690 17.790 19.700 18.000 ;
        RECT 19.850 17.970 20.130 18.260 ;
        RECT 19.870 17.950 20.130 17.970 ;
        RECT 18.550 17.700 19.700 17.790 ;
        RECT 15.330 17.560 19.700 17.700 ;
        RECT 16.320 17.540 19.700 17.560 ;
        RECT 14.250 16.690 16.370 16.960 ;
        RECT 14.250 14.860 14.600 16.690 ;
        RECT 14.850 15.860 15.170 16.190 ;
        RECT 15.330 16.160 16.360 16.690 ;
        RECT 17.090 16.190 17.820 17.540 ;
        RECT 20.380 16.890 21.320 18.720 ;
        RECT 21.570 18.260 21.830 18.290 ;
        RECT 21.570 17.970 21.850 18.260 ;
        RECT 22.010 18.170 23.010 18.720 ;
        RECT 23.880 18.290 24.610 19.640 ;
        RECT 27.100 19.060 27.450 20.890 ;
        RECT 25.330 18.790 27.450 19.060 ;
        RECT 22.010 18.000 23.010 18.010 ;
        RECT 21.570 17.950 21.830 17.970 ;
        RECT 22.000 17.790 23.010 18.000 ;
        RECT 23.150 17.960 25.180 18.290 ;
        RECT 25.340 18.260 26.370 18.790 ;
        RECT 25.355 18.230 26.355 18.260 ;
        RECT 25.355 18.000 26.355 18.020 ;
        RECT 22.000 17.700 23.150 17.790 ;
        RECT 25.330 17.700 26.370 18.000 ;
        RECT 26.530 17.960 26.850 18.290 ;
        RECT 22.000 17.560 26.370 17.700 ;
        RECT 22.000 17.540 25.380 17.560 ;
        RECT 18.690 16.620 23.010 16.890 ;
        RECT 15.345 16.130 16.345 16.160 ;
        RECT 15.345 15.900 16.345 15.920 ;
        RECT 15.330 15.600 16.370 15.900 ;
        RECT 16.520 15.860 18.550 16.190 ;
        RECT 18.690 16.070 19.690 16.620 ;
        RECT 19.870 16.160 20.130 16.190 ;
        RECT 18.690 15.900 19.690 15.910 ;
        RECT 18.690 15.690 19.700 15.900 ;
        RECT 19.850 15.870 20.130 16.160 ;
        RECT 19.870 15.850 20.130 15.870 ;
        RECT 18.550 15.600 19.700 15.690 ;
        RECT 15.330 15.460 19.700 15.600 ;
        RECT 16.320 15.440 19.700 15.460 ;
        RECT 14.250 14.590 16.370 14.860 ;
        RECT 14.250 12.760 14.600 14.590 ;
        RECT 14.850 13.760 15.170 14.090 ;
        RECT 15.330 14.060 16.360 14.590 ;
        RECT 17.090 14.090 17.820 15.440 ;
        RECT 20.380 14.790 21.320 16.620 ;
        RECT 21.570 16.160 21.830 16.190 ;
        RECT 21.570 15.870 21.850 16.160 ;
        RECT 22.010 16.070 23.010 16.620 ;
        RECT 23.880 16.190 24.610 17.540 ;
        RECT 27.100 16.960 27.450 18.790 ;
        RECT 25.330 16.690 27.450 16.960 ;
        RECT 22.010 15.900 23.010 15.910 ;
        RECT 21.570 15.850 21.830 15.870 ;
        RECT 22.000 15.690 23.010 15.900 ;
        RECT 23.150 15.860 25.180 16.190 ;
        RECT 25.340 16.160 26.370 16.690 ;
        RECT 25.355 16.130 26.355 16.160 ;
        RECT 25.355 15.900 26.355 15.920 ;
        RECT 22.000 15.600 23.150 15.690 ;
        RECT 25.330 15.600 26.370 15.900 ;
        RECT 26.530 15.860 26.850 16.190 ;
        RECT 22.000 15.460 26.370 15.600 ;
        RECT 22.000 15.440 25.380 15.460 ;
        RECT 18.690 14.520 23.010 14.790 ;
        RECT 15.345 14.030 16.345 14.060 ;
        RECT 15.345 13.800 16.345 13.820 ;
        RECT 15.330 13.500 16.370 13.800 ;
        RECT 16.520 13.760 18.550 14.090 ;
        RECT 18.690 13.970 19.690 14.520 ;
        RECT 19.870 14.060 20.130 14.090 ;
        RECT 18.690 13.800 19.690 13.810 ;
        RECT 18.690 13.590 19.700 13.800 ;
        RECT 19.850 13.770 20.130 14.060 ;
        RECT 19.870 13.750 20.130 13.770 ;
        RECT 18.550 13.500 19.700 13.590 ;
        RECT 15.330 13.360 19.700 13.500 ;
        RECT 16.320 13.340 19.700 13.360 ;
        RECT 14.250 12.490 16.370 12.760 ;
        RECT 14.250 11.030 14.600 12.490 ;
        RECT 14.850 11.660 15.170 11.990 ;
        RECT 15.330 11.960 16.360 12.490 ;
        RECT 17.090 11.990 17.820 13.340 ;
        RECT 20.380 12.690 21.320 14.520 ;
        RECT 21.570 14.060 21.830 14.090 ;
        RECT 21.570 13.770 21.850 14.060 ;
        RECT 22.010 13.970 23.010 14.520 ;
        RECT 23.880 14.090 24.610 15.440 ;
        RECT 27.100 14.860 27.450 16.690 ;
        RECT 25.330 14.590 27.450 14.860 ;
        RECT 22.010 13.800 23.010 13.810 ;
        RECT 21.570 13.750 21.830 13.770 ;
        RECT 22.000 13.590 23.010 13.800 ;
        RECT 23.150 13.760 25.180 14.090 ;
        RECT 25.340 14.060 26.370 14.590 ;
        RECT 25.355 14.030 26.355 14.060 ;
        RECT 25.355 13.800 26.355 13.820 ;
        RECT 22.000 13.500 23.150 13.590 ;
        RECT 25.330 13.500 26.370 13.800 ;
        RECT 26.530 13.760 26.850 14.090 ;
        RECT 22.000 13.360 26.370 13.500 ;
        RECT 22.000 13.340 25.380 13.360 ;
        RECT 18.690 12.420 23.010 12.690 ;
        RECT 15.345 11.930 16.345 11.960 ;
        RECT 15.345 11.700 16.345 11.720 ;
        RECT 15.330 11.400 16.370 11.700 ;
        RECT 16.520 11.660 18.550 11.990 ;
        RECT 18.690 11.870 19.690 12.420 ;
        RECT 19.870 11.960 20.130 11.990 ;
        RECT 18.690 11.700 19.690 11.710 ;
        RECT 18.690 11.490 19.700 11.700 ;
        RECT 19.850 11.670 20.130 11.960 ;
        RECT 19.870 11.650 20.130 11.670 ;
        RECT 18.550 11.400 19.700 11.490 ;
        RECT 15.330 11.260 19.700 11.400 ;
        RECT 16.320 11.240 19.700 11.260 ;
        RECT 14.240 8.835 14.600 11.030 ;
        RECT 17.090 10.760 17.820 11.240 ;
        RECT 20.380 10.760 21.320 12.420 ;
        RECT 21.570 11.960 21.830 11.990 ;
        RECT 21.570 11.670 21.850 11.960 ;
        RECT 22.010 11.870 23.010 12.420 ;
        RECT 23.880 11.990 24.610 13.340 ;
        RECT 27.100 12.760 27.450 14.590 ;
        RECT 25.330 12.490 27.450 12.760 ;
        RECT 22.010 11.700 23.010 11.710 ;
        RECT 21.570 11.650 21.830 11.670 ;
        RECT 22.000 11.490 23.010 11.700 ;
        RECT 23.150 11.660 25.180 11.990 ;
        RECT 25.340 11.960 26.370 12.490 ;
        RECT 25.355 11.930 26.355 11.960 ;
        RECT 25.355 11.700 26.355 11.720 ;
        RECT 22.000 11.400 23.150 11.490 ;
        RECT 25.330 11.400 26.370 11.700 ;
        RECT 26.530 11.660 26.850 11.990 ;
        RECT 22.000 11.260 26.370 11.400 ;
        RECT 22.000 11.240 25.380 11.260 ;
        RECT 23.880 10.760 24.610 11.240 ;
        RECT 27.100 10.990 27.450 12.490 ;
        RECT 20.380 10.320 21.310 10.760 ;
        RECT 20.380 9.390 21.340 10.320 ;
        RECT 27.090 8.835 27.460 10.990 ;
        RECT 12.645 8.465 27.460 8.835 ;
      LAYER via ;
        RECT 17.170 219.550 17.700 220.620 ;
        RECT 23.960 219.730 24.490 220.680 ;
        RECT 17.140 10.890 17.770 11.300 ;
        RECT 23.950 10.890 24.510 11.320 ;
        RECT 20.520 9.390 21.310 10.320 ;
        RECT 12.675 8.465 13.045 8.835 ;
      LAYER met2 ;
        RECT 17.090 11.390 17.830 220.700 ;
        RECT 23.880 11.400 24.610 220.760 ;
        RECT 17.080 10.760 17.830 11.390 ;
        RECT 17.080 9.890 17.820 10.760 ;
        RECT 20.520 10.320 21.310 10.350 ;
        RECT 12.675 8.835 13.045 8.865 ;
        RECT 12.630 8.465 13.090 8.835 ;
        RECT 12.675 8.435 13.045 8.465 ;
        RECT 17.100 4.820 17.805 9.890 ;
        RECT 20.475 9.390 21.355 10.320 ;
        RECT 20.520 9.360 21.310 9.390 ;
        RECT 23.870 6.220 24.610 11.400 ;
        RECT 23.870 5.500 154.245 6.220 ;
        RECT 23.870 5.490 24.610 5.500 ;
        RECT 17.100 4.125 120.370 4.820 ;
        RECT 17.100 4.120 17.805 4.125 ;
      LAYER via2 ;
        RECT 12.675 8.465 13.045 8.835 ;
        RECT 20.520 9.390 21.310 10.320 ;
        RECT 153.480 5.500 154.200 6.220 ;
        RECT 119.630 4.125 120.325 4.820 ;
      LAYER met3 ;
        RECT 20.495 9.365 21.365 10.345 ;
        RECT 12.580 8.290 13.160 8.940 ;
        RECT 153.455 5.475 154.255 6.245 ;
        RECT 119.605 4.100 120.380 4.845 ;
      LAYER via3 ;
        RECT 20.545 9.365 21.335 10.345 ;
        RECT 12.650 8.440 13.020 8.860 ;
        RECT 153.505 5.475 154.225 6.245 ;
        RECT 119.655 4.100 120.350 4.845 ;
      LAYER met4 ;
        RECT 3.990 223.080 4.290 224.760 ;
        RECT 7.670 223.080 7.970 224.760 ;
        RECT 11.350 223.080 11.650 224.760 ;
        RECT 15.030 223.080 15.330 224.760 ;
        RECT 18.710 223.080 19.010 224.760 ;
        RECT 22.390 223.080 22.690 224.760 ;
        RECT 26.070 223.080 26.370 224.760 ;
        RECT 29.750 223.080 30.050 224.760 ;
        RECT 33.430 223.080 33.730 224.760 ;
        RECT 37.110 223.080 37.410 224.760 ;
        RECT 40.790 223.080 41.090 224.760 ;
        RECT 44.470 223.080 44.770 224.760 ;
        RECT 48.150 223.080 48.450 224.760 ;
        RECT 51.830 223.080 52.130 224.760 ;
        RECT 55.510 223.080 55.810 224.760 ;
        RECT 59.190 223.080 59.490 224.760 ;
        RECT 62.870 223.080 63.170 224.760 ;
        RECT 66.550 223.080 66.850 224.760 ;
        RECT 70.230 223.080 70.530 224.760 ;
        RECT 73.910 223.080 74.210 224.760 ;
        RECT 77.590 223.080 77.890 224.760 ;
        RECT 81.270 223.080 81.570 224.760 ;
        RECT 84.950 223.080 85.250 224.760 ;
        RECT 88.630 223.080 88.930 224.760 ;
        RECT 0.860 221.490 158.950 223.080 ;
        RECT 49.000 220.760 50.500 221.490 ;
        RECT 20.540 10.250 21.340 10.350 ;
        RECT 20.540 9.460 49.000 10.250 ;
        RECT 20.540 9.360 21.340 9.460 ;
        RECT 2.500 8.850 6.890 8.890 ;
        RECT 2.500 8.835 7.960 8.850 ;
        RECT 12.645 8.835 13.025 8.865 ;
        RECT 2.500 8.465 13.025 8.835 ;
        RECT 2.500 8.455 7.960 8.465 ;
        RECT 2.500 8.415 6.890 8.455 ;
        RECT 12.645 8.435 13.025 8.465 ;
        RECT 153.500 6.220 154.230 6.250 ;
        RECT 153.500 5.500 157.040 6.220 ;
        RECT 153.500 5.470 154.230 5.500 ;
        RECT 119.650 4.820 120.355 4.850 ;
        RECT 119.650 4.125 135.105 4.820 ;
        RECT 119.650 4.095 120.355 4.125 ;
        RECT 134.410 1.000 135.105 4.125 ;
        RECT 156.320 1.000 157.040 5.500 ;
        RECT 156.320 0.560 156.410 1.000 ;
  END
END tt_um_devinatkin_dual_oscillator
END LIBRARY

