magic
tech sky130A
magscale 1 2
timestamp 1716415172
<< error_p >>
rect -108 533 -96 545
rect -62 533 62 545
rect 96 533 108 545
rect -133 511 -108 533
rect -96 525 -25 533
rect -62 511 -25 525
rect 25 511 133 533
rect -133 507 -96 511
rect -62 507 133 511
rect -133 501 133 507
rect -162 499 162 501
rect -210 388 -201 499
rect -96 447 -62 478
rect -50 447 50 499
rect 62 447 96 478
rect 108 447 126 477
rect -180 441 -108 447
rect -96 441 22 447
rect 50 441 180 447
rect -180 431 22 441
rect -183 397 -176 404
rect -134 397 -129 431
rect -113 421 -108 431
rect -113 397 -108 407
rect -96 397 -49 431
rect -45 397 22 431
rect -183 388 22 397
rect -210 384 22 388
rect 35 431 180 441
rect 35 397 45 431
rect 62 397 113 431
rect 129 397 134 431
rect 176 397 183 404
rect 35 388 183 397
rect 35 387 209 388
rect -221 350 22 384
rect 50 350 209 387
rect -210 -350 -142 350
rect -134 324 -129 350
rect -109 349 -108 350
rect -96 349 -95 350
rect -63 349 -62 350
rect 62 349 63 350
rect 95 349 96 350
rect 108 349 109 350
rect -28 338 28 349
rect -17 -278 -6 338
rect -129 -324 -6 -278
rect -134 -327 -6 -324
rect 17 -278 28 338
rect 129 324 134 350
rect 142 325 209 350
rect 17 -324 129 -278
rect 17 -327 134 -324
rect -134 -350 134 -327
rect 142 -325 175 325
rect 176 -325 209 325
rect 142 -350 209 -325
rect 210 -350 221 384
rect -210 -351 -107 -350
rect -97 -351 22 -350
rect -210 -387 -108 -351
rect -96 -387 22 -351
rect 50 -387 209 -350
rect -210 -388 22 -387
rect -210 -499 -201 -388
rect -180 -397 22 -388
rect -134 -431 -129 -397
rect -113 -407 -108 -397
rect -113 -431 -108 -421
rect -96 -431 -49 -397
rect -45 -431 22 -397
rect -180 -441 22 -431
rect 35 -388 209 -387
rect 35 -397 180 -388
rect 35 -431 45 -397
rect 62 -431 113 -397
rect 129 -431 134 -397
rect 35 -441 180 -431
rect -180 -447 -108 -441
rect -107 -447 22 -441
rect 50 -447 180 -441
rect -50 -448 -49 -447
rect 49 -448 50 -447
rect -108 -499 -96 -487
rect -62 -499 62 -487
rect 96 -499 108 -487
rect 255 -499 264 499
rect -133 -521 -108 -499
rect -96 -507 -25 -499
rect -62 -521 -25 -507
rect 25 -521 133 -499
rect -133 -525 -96 -521
rect -62 -525 133 -521
rect -133 -533 133 -525
<< nwell >>
rect -246 569 246 969
rect -325 -569 325 569
rect -246 -969 246 -569
<< pmos >>
rect -108 431 -96 447
rect -62 431 -50 447
rect 50 431 62 447
rect 96 431 108 447
rect -108 350 -96 397
rect -62 350 -50 397
rect 50 350 62 397
rect 96 350 108 397
rect -108 -397 -96 -350
rect -62 -397 -50 -350
rect 50 -397 62 -350
rect 96 -397 108 -350
rect -108 -447 -96 -431
rect -62 -447 -50 -431
rect 50 -447 62 -431
rect 96 -447 108 -431
<< pmoslvt >>
rect -50 533 50 750
rect -50 431 50 499
rect -45 397 45 431
rect -50 350 50 397
rect -129 338 129 350
rect -129 -338 -17 338
rect 17 -338 129 338
rect -129 -350 129 -338
rect -50 -397 50 -350
rect -45 -431 45 -397
rect -50 -499 50 -431
rect -50 -750 50 -533
<< pdiff >>
rect -108 738 -50 750
rect -108 533 -96 738
rect -62 533 -50 738
rect 50 738 108 750
rect 50 533 62 738
rect 96 533 108 738
rect -108 447 -96 499
rect -62 447 -50 499
rect 50 447 62 499
rect 96 447 108 499
rect -187 338 -129 350
rect 129 338 187 350
rect -187 -338 -175 338
rect -141 -338 -129 338
rect 129 -338 141 338
rect 175 -338 187 338
rect -187 -350 -129 -338
rect 129 -350 187 -338
rect -108 -499 -96 -447
rect -62 -499 -50 -447
rect 50 -499 62 -447
rect 96 -499 108 -447
rect -108 -738 -96 -533
rect -62 -738 -50 -533
rect -108 -750 -50 -738
rect 50 -738 62 -533
rect 96 -738 108 -533
rect 50 -750 108 -738
<< pdiffc >>
rect -96 533 -62 738
rect 62 533 96 738
rect -96 447 -62 499
rect 62 447 96 499
rect -175 -338 -141 338
rect -17 -338 17 338
rect 141 -338 175 338
rect -96 -499 -62 -447
rect 62 -499 96 -447
rect -96 -738 -62 -533
rect 62 -738 96 -533
<< nsubdiff >>
rect -210 899 -114 933
rect 114 899 210 933
rect -210 837 -176 899
rect 176 837 210 899
rect -289 499 -210 533
rect 210 499 289 533
rect -289 437 -255 499
rect -289 -499 -255 -437
rect 255 437 289 499
rect 255 -499 289 -437
rect -289 -533 -210 -499
rect 210 -533 289 -499
rect -210 -899 -176 -837
rect 176 -899 210 -837
rect -210 -933 -114 -899
rect 114 -933 210 -899
<< nsubdiffcont >>
rect -114 899 114 933
rect -210 533 -176 837
rect 176 533 210 837
rect -210 499 210 533
rect -289 -437 -255 437
rect -210 350 -176 499
rect 176 350 210 499
rect -210 -350 -187 350
rect 187 -350 210 350
rect -210 -499 -176 -350
rect 176 -499 210 -350
rect 255 -437 289 437
rect -210 -533 210 -499
rect -210 -837 -176 -533
rect 176 -837 210 -533
rect -114 -933 114 -899
<< poly >>
rect -50 831 50 847
rect -50 797 -34 831
rect 34 797 50 831
rect -50 750 50 797
rect -129 431 -108 447
rect -96 431 -62 447
rect 62 431 96 447
rect 108 431 129 447
rect -129 397 -113 431
rect 113 397 129 431
rect -129 350 -108 397
rect -96 350 -62 397
rect 62 350 96 397
rect 108 350 129 397
rect -129 -397 -108 -350
rect -96 -397 -62 -350
rect 62 -397 96 -350
rect 108 -397 129 -350
rect -129 -431 -113 -397
rect 113 -431 129 -397
rect -129 -447 -108 -431
rect -96 -447 -62 -431
rect 62 -447 96 -431
rect 108 -447 129 -431
rect -50 -797 50 -750
rect -50 -831 -34 -797
rect 34 -831 50 -797
rect -50 -847 50 -831
<< polycont >>
rect -34 797 34 831
rect -113 397 -45 431
rect 45 397 113 431
rect -113 -431 -45 -397
rect 45 -431 113 -397
rect -34 -831 34 -797
<< locali >>
rect -210 899 -114 933
rect 114 899 210 933
rect -210 837 -176 899
rect 176 837 210 899
rect -50 797 -34 831
rect 34 797 50 831
rect -96 738 -62 754
rect 62 738 96 754
rect -289 499 -210 533
rect 210 499 289 533
rect -289 437 -255 499
rect -289 -499 -255 -437
rect -129 397 -113 431
rect -45 397 -29 431
rect 29 397 45 431
rect 113 397 129 431
rect -187 -350 -176 350
rect -175 338 -141 354
rect -175 -354 -141 -338
rect -17 338 17 354
rect -17 -354 17 -338
rect 141 338 175 354
rect 141 -354 175 -338
rect 176 -350 187 350
rect -129 -431 -113 -397
rect -45 -431 -29 -397
rect 29 -431 45 -397
rect 113 -431 129 -397
rect 255 437 289 499
rect 255 -499 289 -437
rect -289 -533 -210 -499
rect 210 -533 289 -499
rect -96 -754 -62 -738
rect 62 -754 96 -738
rect -50 -831 -34 -797
rect 34 -831 50 -797
rect -210 -899 -176 -837
rect 176 -899 210 -837
rect -210 -933 -114 -899
rect 114 -933 210 -899
<< viali >>
rect -34 797 34 831
rect -96 533 -62 738
rect 62 533 96 738
rect -96 499 -62 533
rect 62 499 96 533
rect -96 447 -62 499
rect -96 431 -62 447
rect 62 447 96 499
rect 62 431 96 447
rect -113 397 -45 431
rect 45 397 113 431
rect -175 -338 -141 338
rect -96 -397 -62 397
rect -17 -338 17 338
rect 62 -397 96 397
rect 141 -338 175 338
rect -113 -431 -45 -397
rect 45 -431 113 -397
rect -96 -447 -62 -431
rect -96 -499 -62 -447
rect 62 -447 96 -431
rect 62 -499 96 -447
rect -96 -533 -62 -499
rect 62 -533 96 -499
rect -96 -738 -62 -533
rect 62 -738 96 -533
rect -34 -831 34 -797
<< metal1 >>
rect -46 831 46 837
rect -46 797 -34 831
rect 34 797 46 831
rect -46 791 46 797
rect -102 738 -56 750
rect -102 437 -96 738
rect -125 431 -96 437
rect -62 437 -56 738
rect 56 738 102 750
rect 56 437 62 738
rect -62 431 -33 437
rect -125 397 -113 431
rect -45 397 -33 431
rect -125 391 -96 397
rect -181 338 -135 350
rect -181 -338 -175 338
rect -141 -338 -135 338
rect -181 -350 -135 -338
rect -102 -391 -96 391
rect -125 -397 -96 -391
rect -62 391 -33 397
rect 33 431 62 437
rect 96 437 102 738
rect 96 431 125 437
rect 33 397 45 431
rect 113 397 125 431
rect 33 391 62 397
rect -62 -391 -56 391
rect -23 338 23 350
rect -23 -338 -17 338
rect 17 -338 23 338
rect -23 -350 23 -338
rect 56 -391 62 391
rect -62 -397 -33 -391
rect -125 -431 -113 -397
rect -45 -431 -33 -397
rect -125 -437 -96 -431
rect -102 -738 -96 -437
rect -62 -437 -33 -431
rect 33 -397 62 -391
rect 96 391 125 397
rect 96 -391 102 391
rect 135 338 181 350
rect 135 -338 141 338
rect 175 -338 181 338
rect 135 -350 181 -338
rect 96 -397 125 -391
rect 33 -431 45 -397
rect 113 -431 125 -397
rect 33 -437 62 -431
rect -62 -738 -56 -437
rect -102 -750 -56 -738
rect 56 -738 62 -437
rect 96 -437 125 -431
rect 96 -738 102 -437
rect 56 -750 102 -738
rect -46 -797 46 -791
rect -46 -831 -34 -797
rect 34 -831 46 -797
rect -46 -837 46 -831
<< properties >>
string FIXED_BBOX -272 -516 272 516
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 3.5 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
