magic
tech sky130A
magscale 1 2
timestamp 1716521300
<< error_p >>
rect -34 546 34 547
rect -50 -500 50 -499
<< nwell >>
rect -144 -600 144 600
<< pmoslvt >>
rect -50 -500 50 500
<< pdiff >>
rect -108 488 -50 500
rect -108 -488 -96 488
rect -62 -488 -50 488
rect -108 -500 -50 -488
rect 50 488 108 500
rect 50 -488 62 488
rect 96 -488 108 488
rect 50 -500 108 -488
<< pdiffc >>
rect -96 -488 -62 488
rect 62 -488 96 488
<< poly >>
rect -50 580 50 596
rect -50 546 -34 580
rect 34 546 50 580
rect -50 500 50 546
rect -50 -546 50 -500
rect -50 -580 -34 -546
rect 34 -580 50 -546
rect -50 -596 50 -580
<< polycont >>
rect -34 546 34 580
rect -34 -580 34 -546
<< locali >>
rect -50 546 -34 580
rect 34 546 50 580
rect -96 488 -62 504
rect -96 -504 -62 -488
rect 62 488 96 504
rect 62 -504 96 -488
rect -50 -580 -34 -546
rect 34 -580 50 -546
<< viali >>
rect -34 546 34 580
rect -96 -488 -62 488
rect 62 -488 96 488
rect -34 -580 34 -546
<< metal1 >>
rect -46 580 46 586
rect -46 546 -34 580
rect 34 546 46 580
rect -46 540 46 546
rect -102 488 -56 500
rect -102 -488 -96 488
rect -62 -488 -56 488
rect -102 -500 -56 -488
rect 56 488 102 500
rect 56 -488 62 488
rect 96 -488 102 488
rect 56 -500 102 -488
rect -46 -546 46 -540
rect -46 -580 -34 -546
rect 34 -580 46 -546
rect -46 -586 46 -580
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
