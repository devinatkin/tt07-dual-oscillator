magic
tech sky130A
magscale 1 2
timestamp 1716524512
<< pwell >>
rect 1090 -540 1416 -430
<< metal1 >>
rect 430 6048 554 6238
rect 8005 6126 8186 6204
rect 439 5375 545 6048
rect 442 2074 542 5375
rect 443 165 542 2074
rect 8005 409 8083 6126
rect 8241 4506 8319 4512
rect 8319 4428 8650 4506
rect 8241 4422 8319 4428
rect 12914 3242 13300 3272
rect 12914 2936 12976 3242
rect 13258 3136 13300 3242
rect 13258 2948 15962 3136
rect 13258 2936 13300 2948
rect 12914 2892 13300 2936
rect 8005 325 8083 331
rect -151 35 543 165
rect 15774 152 15962 2948
rect 820 52 1056 84
rect -151 -48 -21 35
rect -266 -168 94 -48
rect 820 -116 846 52
rect 1032 -116 1056 52
rect 820 -146 1056 -116
rect 9260 -70 9532 60
rect 15774 -29 20555 152
rect 15774 -33 15962 -29
rect -758 -742 94 -168
rect 9260 -160 9276 -70
rect 9514 -160 9532 -70
rect 9260 -176 9532 -160
rect 19162 -207 19358 -206
rect 496 -430 15508 -374
rect 18894 -403 18900 -207
rect 19096 -403 19358 -207
rect 404 -458 15508 -430
rect 404 -528 1164 -458
rect 1292 -484 15508 -458
rect 1292 -528 1416 -484
rect 404 -538 1416 -528
rect 1090 -540 1416 -538
rect -266 -1896 94 -742
rect 19162 -1120 19358 -403
rect 18346 -1316 19358 -1120
rect 20374 -1752 20555 -29
rect -266 -1904 764 -1896
rect -266 -2246 1350 -1904
rect 20374 -1933 26896 -1752
rect 7791 -2097 7797 -2019
rect 7875 -2097 7881 -2019
rect -266 -2256 764 -2246
rect 26715 -2576 26896 -1933
rect 26718 -2862 26892 -2576
rect 26296 -3064 26892 -2862
rect -1384 -3634 -1236 -3610
rect -534 -3634 622 -3610
rect -1384 -3724 622 -3634
rect 1098 -3624 1326 -3612
rect 1098 -3700 1164 -3624
rect 1296 -3700 1326 -3624
rect 1098 -3716 1326 -3700
<< via1 >>
rect 8241 4428 8319 4506
rect 12976 2936 13258 3242
rect 8005 331 8083 409
rect 846 -116 1032 52
rect 9276 -160 9514 -70
rect 18900 -403 19096 -207
rect 1164 -528 1292 -458
rect 7797 -2097 7875 -2019
rect -936 -3572 -618 -3166
rect 1164 -3700 1296 -3624
<< metal2 >>
rect 964 3332 1022 4454
rect 8235 4428 8241 4506
rect 8319 4428 8325 4506
rect 284 3202 544 3240
rect 284 2970 318 3202
rect 494 2970 544 3202
rect 284 2938 544 2970
rect 300 532 497 2938
rect 964 1694 1024 3332
rect 894 1664 1122 1694
rect 894 1466 912 1664
rect 1088 1466 1122 1664
rect 8241 1683 8319 4428
rect 12914 3242 13300 3272
rect 12914 2936 12976 3242
rect 13258 2936 13300 3242
rect 12914 2892 13300 2936
rect 8241 1596 8319 1605
rect 894 1448 1122 1466
rect 300 225 496 532
rect 7999 331 8005 409
rect 8083 331 8089 409
rect 296 39 305 225
rect 491 39 500 225
rect 804 52 1058 84
rect 300 34 496 39
rect 804 -24 846 52
rect -994 -116 846 -24
rect 1032 -116 1058 52
rect -994 -146 1058 -116
rect -988 -742 -558 -146
rect 8005 -273 8083 331
rect 9260 -70 9532 -60
rect 9260 -160 9276 -70
rect 9514 -160 9532 -70
rect 9260 -176 9532 -160
rect 7797 -351 8083 -273
rect 18868 -207 19124 -176
rect 1144 -458 1308 -446
rect 1144 -528 1164 -458
rect 1292 -528 1308 -458
rect -988 -1422 -806 -742
rect -988 -3166 -558 -1422
rect -988 -3572 -936 -3166
rect -618 -3572 -558 -3166
rect -988 -3592 -558 -3572
rect 1144 -3624 1308 -528
rect 7797 -2019 7875 -351
rect 18868 -403 18900 -207
rect 19096 -403 19124 -207
rect 18868 -434 19124 -403
rect 7797 -2103 7875 -2097
rect 1144 -3700 1164 -3624
rect 1296 -3700 1308 -3624
rect 1144 -3706 1308 -3700
<< via2 >>
rect 318 2970 494 3202
rect 912 1466 1088 1664
rect 12976 2936 13258 3242
rect 8241 1605 8319 1683
rect 305 39 491 225
rect 850 -114 1024 18
rect 9276 -160 9514 -70
rect 18900 -403 19096 -207
<< metal3 >>
rect 12914 3264 13300 3272
rect 10294 3242 13300 3264
rect 284 3202 544 3240
rect 284 2970 318 3202
rect 494 3098 544 3202
rect 494 2994 2800 3098
rect 494 2970 544 2994
rect 10294 2982 12976 3242
rect 284 2938 544 2970
rect 12914 2936 12976 2982
rect 13258 2936 13300 3242
rect 12914 2892 13300 2936
rect 6882 1716 7950 1720
rect 786 1664 7950 1716
rect 786 1466 912 1664
rect 1088 1468 7950 1664
rect 8236 1683 8324 1688
rect 14724 1683 15792 1720
rect 8236 1605 8241 1683
rect 8319 1605 15792 1683
rect 8236 1600 8324 1605
rect 14724 1468 15792 1605
rect 1088 1466 7438 1468
rect 786 1458 7438 1466
rect 786 1434 4638 1458
rect 5102 1434 7438 1458
rect 300 225 496 230
rect 300 39 305 225
rect 491 39 496 225
rect 300 -208 496 39
rect 800 18 1104 40
rect 800 -114 850 18
rect 1024 14 1104 18
rect 1024 -114 1118 14
rect 800 -144 1118 -114
rect 300 -402 301 -208
rect 495 -402 496 -208
rect 300 -403 496 -402
rect 908 -198 1118 -144
rect 9258 -70 9532 -44
rect 9258 -160 9276 -70
rect 9514 -160 9532 -70
rect 908 -342 1300 -198
rect 9258 -342 9532 -160
rect 18868 -202 19124 -176
rect 301 -408 495 -403
rect 908 -534 10032 -342
rect 18868 -408 18895 -202
rect 19101 -408 19124 -202
rect 18868 -434 19124 -408
<< via3 >>
rect 301 -402 495 -208
rect 18895 -207 19101 -202
rect 18895 -403 18900 -207
rect 18900 -403 19096 -207
rect 19096 -403 19101 -207
rect 18895 -408 19101 -403
<< metal4 >>
rect 18894 -202 19102 -201
rect 18894 -207 18895 -202
rect 300 -208 18895 -207
rect 300 -402 301 -208
rect 495 -402 18895 -208
rect 300 -403 18895 -402
rect 18894 -408 18895 -403
rect 19101 -408 19102 -202
rect 18894 -409 19102 -408
use current_source  current_source_0
timestamp 1716523272
transform 1 0 -1330 0 1 -4270
box -54 544 936 8966
use opamp_1  opamp_1_0
timestamp 1716526700
transform 1 0 6896 0 1 2202
box 1092 -2630 8676 5872
use opamp_1  opamp_1_1
timestamp 1716526700
transform 1 0 -688 0 1 2202
box 1092 -2630 8676 5872
use oscillator_20MHZ  oscillator_20MHZ_0
timestamp 1716523272
transform 1 0 404 0 1 -3721
box 0 -1 26159 1646
use oscillator_21MHZ  oscillator_21MHZ_0
timestamp 1716523272
transform 1 0 404 0 -1 -431
box 0 -1 18074 1645
<< labels >>
flabel metal1 428 -2228 1106 -1930 0 FreeSans 1600 0 0 0 VCC
port 0 nsew
flabel metal1 1098 -3716 1326 -3612 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal3 6882 1468 7950 1720 0 FreeSans 480 0 0 0 OUTB
port 6 nsew
flabel metal3 14724 1468 15792 1720 0 FreeSans 480 0 0 0 OUTA
port 5 nsew
<< end >>
