magic
tech sky130A
magscale 1 2
timestamp 1716849570
<< metal1 >>
rect 19306 30088 19818 30158
rect 19306 29660 19382 30088
rect 19734 29660 19818 30088
rect 19306 29596 19818 29660
rect 17536 29318 17938 29372
rect 17536 28646 17584 29318
rect 17726 28646 17938 29318
rect 17536 28604 17938 28646
<< via1 >>
rect 19382 29660 19734 30088
rect 17584 28646 17726 29318
<< metal2 >>
rect 19306 30088 19818 30158
rect 19306 29660 19382 30088
rect 19734 29660 19818 30088
rect 19306 29596 19818 29660
rect 17538 29318 17784 29378
rect 17538 28646 17584 29318
rect 17726 28646 17784 29318
rect 17538 28610 17784 28646
<< via2 >>
rect 19384 29662 19734 30088
rect 17584 28646 17726 29318
<< metal3 >>
rect 19306 30134 19818 30158
rect 176 30098 19818 30134
rect 176 29672 242 30098
rect 466 30088 19818 30098
rect 466 29672 19384 30088
rect 176 29662 19384 29672
rect 19734 29662 19818 30088
rect 176 29638 19818 29662
rect 500 29634 19818 29638
rect 19306 29596 19818 29634
rect 17538 29318 17784 29378
rect 17538 29264 17584 29318
rect 9802 29218 17584 29264
rect 9802 28718 9840 29218
rect 10048 28718 17584 29218
rect 9802 28692 17584 28718
rect 17538 28646 17584 28692
rect 17726 28646 17784 29318
rect 17538 28610 17784 28646
rect 23064 21763 24018 21836
rect 23064 21644 25166 21763
rect 23784 21624 25166 21644
rect 23784 21529 28807 21624
rect 25074 21468 28806 21529
rect 26410 21374 28806 21468
rect 23064 13296 23316 14236
rect 23070 1626 23310 13296
rect 26840 2334 27086 2354
rect 28575 2334 28806 21374
rect 26560 2306 28806 2334
rect 26560 2108 26884 2306
rect 27032 2108 28806 2306
rect 26560 2103 28806 2108
rect 26560 2098 28644 2103
rect 26840 2074 27086 2098
rect 31222 1626 31476 1642
rect 23070 1596 31678 1626
rect 23070 1410 31268 1596
rect 31422 1410 31678 1596
rect 23070 1386 31678 1410
rect 31222 1362 31476 1386
<< via3 >>
rect 242 29672 466 30098
rect 9840 28718 10048 29218
rect 26884 2108 27032 2306
rect 31268 1410 31422 1596
<< metal4 >>
rect 798 44644 858 45152
rect 1534 44644 1594 45152
rect 2270 44644 2330 45152
rect 3006 44644 3066 45152
rect 3742 44644 3802 45152
rect 4478 44644 4538 45152
rect 5214 44644 5274 45152
rect 5950 44644 6010 45152
rect 6686 44644 6746 45152
rect 7422 44644 7482 45152
rect 8158 44644 8218 45152
rect 8894 44644 8954 45152
rect 9630 44644 9690 45152
rect 10366 44644 10426 45152
rect 11102 44644 11162 45152
rect 11838 44644 11898 45152
rect 12574 44644 12634 45152
rect 13310 44644 13370 45152
rect 14046 44644 14106 45152
rect 14782 44644 14842 45152
rect 15518 44644 15578 45152
rect 16254 44644 16314 45152
rect 16990 44644 17050 45152
rect 17726 44644 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 594 44324 17918 44644
rect 200 30098 500 44152
rect 200 29672 242 30098
rect 466 29672 500 30098
rect 200 1000 500 29672
rect 9800 29218 10100 44324
rect 9800 28718 9840 29218
rect 10048 28718 10100 29218
rect 9800 1000 10100 28718
rect 26840 2306 27086 2354
rect 26840 2108 26884 2306
rect 27032 2108 27086 2306
rect 26840 2074 27086 2108
rect 26869 499 27044 2074
rect 31222 1596 31476 1642
rect 31222 1410 31268 1596
rect 31422 1410 31476 1596
rect 31222 1362 31476 1410
rect 26871 200 27041 499
rect 31307 200 31426 1362
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 200
use top  top_0 ~/tt07-dual-oscillator/mag
timestamp 1716849570
transform 0 1 21596 -1 0 29776
box -1384 -3733 26896 8074
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 200 1000 500 44152 0 FreeSans 1600 0 0 0 VPWR
port 53 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
