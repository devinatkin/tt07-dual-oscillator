magic
tech sky130A
magscale 1 2
timestamp 1716506148
<< pwell >>
rect -739 -692 739 692
<< psubdiff >>
rect -703 622 -607 656
rect 607 622 703 656
rect -703 560 -669 622
rect 669 560 703 622
rect -703 -622 -669 -560
rect 669 -622 703 -560
rect -703 -656 -607 -622
rect 607 -656 703 -622
<< psubdiffcont >>
rect -607 622 607 656
rect -703 -560 -669 560
rect 669 -560 703 560
rect -607 -656 607 -622
<< xpolycontact >>
rect -573 94 573 526
rect -573 -526 573 -94
<< xpolyres >>
rect -573 -94 573 94
<< locali >>
rect -703 622 -607 656
rect 607 622 703 656
rect -703 560 -669 622
rect 669 560 703 622
rect -703 -622 -669 -560
rect 669 -622 703 -560
rect -703 -656 -607 -622
rect 607 -656 703 -622
<< viali >>
rect -557 111 557 508
rect -557 -508 557 -111
<< metal1 >>
rect -569 508 569 514
rect -569 111 -557 508
rect 557 111 569 508
rect -569 105 569 111
rect -569 -111 569 -105
rect -569 -508 -557 -111
rect 557 -508 569 -111
rect -569 -514 569 -508
<< properties >>
string FIXED_BBOX -686 -639 686 639
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 1.1 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 449.633 dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
