magic
tech sky130A
timestamp 1717178954
<< metal1 >>
rect 183 5383 398 5596
rect 2899 5546 3441 5596
rect 2899 5259 3114 5436
rect 183 5249 3114 5259
rect 183 5190 2912 5249
rect 3104 5190 3114 5249
rect 183 5183 3114 5190
rect 3226 5186 3441 5435
rect 5941 5383 6156 5596
rect 183 4972 398 5183
rect 3226 5182 5267 5186
rect 3254 5181 5267 5182
rect 3254 5129 5221 5181
rect 5260 5129 5267 5181
rect 3254 5125 5267 5129
rect 5319 5161 5373 5169
rect 183 4646 398 4859
rect 2898 4809 3113 5022
rect 184 4400 398 4533
rect 2898 4483 3113 4696
rect 0 4271 398 4400
rect 1004 4360 1337 4361
rect 3254 4360 3322 5125
rect 5319 5124 5328 5161
rect 5363 5150 5373 5161
rect 5363 5125 6249 5150
rect 5363 5124 5373 5125
rect 5319 5114 5373 5124
rect 941 4348 3322 4360
rect 941 4301 953 4348
rect 1067 4301 3322 4348
rect 941 4292 3322 4301
rect 3895 4957 4158 5019
rect 4220 4957 4223 5019
rect 941 4291 1337 4292
rect 42 4162 1487 4220
rect 3895 1076 3957 4957
rect 3653 1075 3957 1076
rect 3469 1058 3957 1075
rect 3469 960 3483 1058
rect 3607 1014 3957 1058
rect 5374 1111 5411 1115
rect 3607 1013 3752 1014
rect 3607 960 3619 1013
rect 3469 949 3619 960
rect 5374 1000 5376 1111
rect 5409 1000 5411 1111
rect 273 213 1275 253
rect 5374 62 5411 1000
rect 3667 43 6890 62
rect -1 1 6890 43
<< via1 >>
rect 2912 5190 3104 5249
rect 5221 5129 5260 5181
rect 5328 5124 5363 5161
rect 953 4301 1067 4348
rect 4158 4957 4220 5019
rect 3483 960 3607 1058
rect 5376 1000 5409 1111
<< metal2 >>
rect 2899 5249 3114 5259
rect 2899 5190 2912 5249
rect 3104 5190 3114 5249
rect 2899 5183 3114 5190
rect 5218 5181 5267 5186
rect 5218 5129 5221 5181
rect 5260 5129 5267 5181
rect 5218 5125 5267 5129
rect 5319 5161 5373 5169
rect 5319 5124 5328 5161
rect 5363 5124 5373 5161
rect 5319 5114 5373 5124
rect 4158 5019 4220 5022
rect 5294 5019 5334 5114
rect 4220 4957 5334 5019
rect 4158 4954 4220 4957
rect 941 4348 1080 4360
rect 941 4301 953 4348
rect 1067 4301 1080 4348
rect 941 4291 1080 4301
rect 941 3042 965 4291
rect 941 3015 1010 3042
rect 982 2934 1010 3015
rect 244 2392 379 2503
rect 274 1020 311 2392
rect 982 2372 1011 2934
rect 982 2338 1122 2372
rect 1072 1709 1122 2338
rect 5369 1111 5413 1115
rect 3469 1058 3619 1075
rect 274 1016 351 1020
rect 274 975 279 1016
rect 342 975 351 1016
rect 274 970 351 975
rect 3469 960 3483 1058
rect 3607 960 3619 1058
rect 5369 1000 5376 1111
rect 5409 1000 5413 1111
rect 5369 996 5413 1000
rect 3469 949 3619 960
<< via2 >>
rect 2912 5190 3104 5249
rect 5223 5132 5256 5178
rect 5328 5124 5363 5161
rect 279 975 342 1016
rect 3483 960 3607 1058
rect 5376 1007 5409 1102
<< metal3 >>
rect 2899 5249 3114 5259
rect 2899 5190 2912 5249
rect 3104 5234 3114 5249
rect 3104 5228 5139 5234
rect 3104 5191 5094 5228
rect 5133 5191 5139 5228
rect 3104 5190 5139 5191
rect 2899 5184 5139 5190
rect 2899 5183 3114 5184
rect 5218 5178 5267 5186
rect 5218 5132 5223 5178
rect 5256 5132 5267 5178
rect 5218 5125 5267 5132
rect 5319 5161 5373 5169
rect 5319 5124 5328 5161
rect 5363 5124 5373 5161
rect 5319 5114 5373 5124
rect 5369 1102 5413 1115
rect 3305 1058 3618 1074
rect 3305 1020 3483 1058
rect 263 1016 3483 1020
rect 263 975 279 1016
rect 342 975 3483 1016
rect 263 970 3483 975
rect 3305 960 3483 970
rect 3607 1020 3618 1058
rect 3607 970 3619 1020
rect 5369 1007 5376 1102
rect 5409 1007 5413 1102
rect 5369 996 5413 1007
rect 3607 960 3618 970
rect 3305 948 3618 960
<< via3 >>
rect 5094 5191 5133 5228
rect 5223 5132 5256 5178
rect 5328 5124 5363 5161
<< metal4 >>
rect 5089 5228 5163 5234
rect 5089 5191 5094 5228
rect 5133 5191 5163 5228
rect 5089 5188 5163 5191
rect 5113 5047 5163 5188
rect 5218 5178 5267 5186
rect 5218 5132 5223 5178
rect 5256 5132 5267 5178
rect 5218 4995 5267 5132
rect 5319 5161 5373 5169
rect 5319 5124 5328 5161
rect 5363 5124 5373 5161
rect 5319 5114 5373 5124
rect 5319 5007 5358 5114
use capacitor_array  capacitor_array_0
timestamp 1717178954
transform -1 0 6666 0 -1 4853
box -248 -210 2818 4670
use opamp_1  opamp_1_0
timestamp 1717178954
transform 1 0 -546 0 1 1315
box 546 -1315 4338 2936
use sky130_fd_pr__res_generic_po_FKS477  sky130_fd_pr__res_generic_po_FKS477_0
timestamp 1717178954
transform 0 -1 1648 1 0 5571
box -108 -1548 108 1548
use sky130_fd_pr__res_generic_po_FKS477  sky130_fd_pr__res_generic_po_FKS477_1
timestamp 1717178954
transform 0 -1 1648 1 0 4508
box -108 -1548 108 1548
use sky130_fd_pr__res_generic_po_FKS477  sky130_fd_pr__res_generic_po_FKS477_2
timestamp 1717178954
transform 0 -1 1648 1 0 4671
box -108 -1548 108 1548
use sky130_fd_pr__res_generic_po_FKS477  sky130_fd_pr__res_generic_po_FKS477_3
timestamp 1717178954
transform 0 -1 1648 1 0 4834
box -108 -1548 108 1548
use sky130_fd_pr__res_generic_po_FKS477  sky130_fd_pr__res_generic_po_FKS477_4
timestamp 1717178954
transform 0 -1 1648 1 0 4997
box -108 -1548 108 1548
use sky130_fd_pr__res_generic_po_FKS477  sky130_fd_pr__res_generic_po_FKS477_5
timestamp 1717178954
transform 0 -1 1648 1 0 5408
box -108 -1548 108 1548
use sky130_fd_pr__res_generic_po_FKS477  sky130_fd_pr__res_generic_po_FKS477_6
timestamp 1717178954
transform 0 -1 4691 1 0 5408
box -108 -1548 108 1548
use sky130_fd_pr__res_generic_po_FKS477  sky130_fd_pr__res_generic_po_FKS477_7
timestamp 1717178954
transform 0 -1 4691 1 0 5571
box -108 -1548 108 1548
<< labels >>
flabel metal1 183 5183 3114 5259 0 FreeSans 800 0 0 0 mid
flabel metal1 0 4271 398 4400 0 FreeSans 800 0 0 0 fil_in
port 1 nsew
flabel metal1 3226 5182 3441 5435 0 FreeSans 800 0 0 0 op_inb
flabel metal1 -1 1 3761 43 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel metal1 42 4162 1487 4220 0 FreeSans 800 0 0 0 VCC
port 3 nsew
flabel metal3 263 970 746 1019 0 FreeSans 800 0 0 0 fil_out
port 4 nsew
flabel metal1 5329 5125 6249 5150 0 FreeSans 800 0 0 0 fil_out
port 5 nsew
flabel metal1 273 213 1275 253 0 FreeSans 800 0 0 0 IBIAS
port 6 nsew
<< end >>
