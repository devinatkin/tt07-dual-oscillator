magic
tech sky130A
magscale 1 2
timestamp 1717178954
<< nwell >>
rect 22578 8482 22974 11902
rect 14980 5040 15368 7290
rect 18276 1636 18992 1916
<< pwell >>
rect 15034 7290 15150 11902
<< metal1 >>
rect 12448 22430 12692 22480
rect 12448 22238 12484 22430
rect 12650 22238 12692 22430
rect 12448 22200 12692 22238
rect 15404 22428 15678 22480
rect 15404 22266 15448 22428
rect 15656 22302 15678 22428
rect 15656 22266 15770 22302
rect 15404 22252 15770 22266
rect 15404 22224 15678 22252
rect 30838 20854 31168 20898
rect -482 20774 176 20802
rect 30838 20800 30894 20854
rect -1260 20566 -866 20608
rect -1260 20206 -1196 20566
rect -920 20440 -866 20566
rect -482 20596 -366 20774
rect 128 20596 176 20774
rect -482 20554 176 20596
rect 27506 20546 30894 20800
rect 30838 20530 30894 20546
rect 31122 20530 31168 20854
rect 30838 20466 31168 20530
rect 28298 20442 28834 20454
rect -920 20324 150 20440
rect 27776 20326 28834 20442
rect -920 20206 -866 20324
rect -1260 20172 -866 20206
rect 28298 17214 28834 20326
rect 28298 16650 29810 17214
rect 28366 13470 29326 16650
rect 20550 13434 20722 13452
rect 7344 13398 7588 13414
rect 7344 13304 7372 13398
rect 7562 13304 7588 13398
rect 7344 13288 7588 13304
rect 20550 13304 20574 13434
rect 20696 13350 20722 13434
rect 20696 13304 20910 13350
rect 20550 13284 20910 13304
rect 28366 13002 28550 13470
rect 29202 13002 29326 13470
rect 28366 12928 29326 13002
rect 29614 13706 30026 13782
rect 29614 12276 29684 13706
rect 29966 12276 30026 13706
rect 29614 12216 30026 12276
rect 28586 12126 29852 12128
rect 13638 12002 14532 12126
rect 27476 12006 29852 12126
rect 27476 12004 28742 12006
rect 25696 11838 29418 11858
rect 188 11822 29418 11838
rect 188 11724 28520 11822
rect 188 11690 4552 11724
rect 4306 11650 4362 11690
rect 11308 11672 13954 11724
rect 16280 11654 19770 11724
rect 25696 11662 28520 11724
rect 29240 11662 29418 11822
rect 29710 11744 29852 12006
rect 30338 11744 30418 12136
rect 30696 11822 31318 11858
rect 30696 11744 30746 11822
rect 29710 11676 30746 11744
rect 25696 11630 29418 11662
rect 29752 11602 30746 11676
rect 30394 11600 30746 11602
rect 30696 11570 30746 11600
rect 31286 11570 31318 11822
rect 30696 11538 31318 11570
rect 3078 7170 3362 7220
rect 3078 6462 3104 7170
rect 3322 6462 3362 7170
rect 5210 6976 5490 7006
rect 5210 6806 5250 6976
rect 5444 6806 5490 6976
rect 5210 6784 5490 6806
rect 27076 6816 27366 6882
rect 14924 6542 15220 6562
rect 14924 6474 14954 6542
rect 3078 6424 3362 6462
rect 14088 6414 14954 6474
rect 15190 6474 15220 6542
rect 15190 6414 15798 6474
rect 14088 6390 15798 6414
rect 27076 6432 27126 6816
rect 27316 6432 27366 6816
rect 27076 6396 27366 6432
rect 14924 6388 15220 6390
rect -432 4940 -146 4972
rect -432 4704 -390 4940
rect -180 4862 -146 4940
rect 30474 4900 30656 4938
rect 30474 4864 30504 4900
rect -180 4704 3188 4862
rect 12024 4708 18588 4858
rect 27274 4720 30504 4864
rect 30474 4716 30504 4720
rect 30624 4716 30656 4900
rect -432 4692 3188 4704
rect -432 4670 -146 4692
rect 30474 4676 30656 4716
rect 6612 3436 7804 3524
rect 9718 3444 11624 3450
rect 7846 3442 11624 3444
rect 7846 3436 13474 3442
rect 5994 3426 13474 3436
rect 14812 3440 16004 3524
rect 14812 3434 20286 3440
rect 22510 3434 23702 3524
rect 14812 3426 24026 3434
rect 5994 3422 24026 3426
rect 5994 3278 24074 3422
rect 5994 3264 18236 3278
rect 5994 3258 9752 3264
rect 5994 3250 7900 3258
rect 11568 3256 18236 3264
rect 13404 3242 18236 3256
rect 13404 3240 15310 3242
rect 18200 3130 18236 3242
rect 18560 3242 24074 3278
rect 18560 3130 18580 3242
rect 20158 3222 24026 3242
rect 18200 3102 18580 3130
rect 24328 2774 24778 2802
rect 24328 2594 24388 2774
rect 23968 2400 24388 2594
rect 24328 2334 24388 2400
rect 24740 2334 24778 2774
rect 24328 2282 24778 2334
rect 3000 1912 3836 1974
rect -1442 1776 -820 1820
rect -1442 1702 -1394 1776
rect -1470 1508 -1394 1702
rect -1442 1446 -1394 1508
rect -862 1702 -820 1776
rect 3000 1702 3078 1912
rect -862 1672 3078 1702
rect 3768 1672 3836 1912
rect 26874 1842 27270 1878
rect -862 1618 3836 1672
rect -862 1508 3532 1618
rect 26874 1602 26916 1842
rect 27242 1602 27270 1842
rect 26874 1564 27270 1602
rect -862 1446 -820 1508
rect 26576 1464 26776 1560
rect 28200 1462 28400 1558
rect -1442 1406 -820 1446
rect 2046 946 2394 988
rect 2046 598 2094 946
rect 2358 860 2394 946
rect 2358 660 3200 860
rect 2358 598 2394 660
rect 2046 558 2394 598
rect 18198 206 18582 238
rect 18198 32 18238 206
rect 18554 32 18582 206
rect 30696 142 31318 170
rect 30696 108 30738 142
rect 18198 0 18582 32
rect 28946 2 30738 108
rect 30696 -20 30738 2
rect 31282 -20 31318 142
rect 30696 -42 31318 -20
<< via1 >>
rect 12484 22238 12650 22430
rect 15448 22266 15656 22428
rect -1196 20206 -920 20566
rect -366 20596 128 20774
rect 30894 20530 31122 20854
rect 29734 19740 29898 20022
rect 7372 13304 7562 13398
rect 20574 13304 20696 13434
rect 28550 13002 29202 13470
rect 29684 12276 29966 13706
rect 28520 11662 29240 11822
rect 30746 11570 31286 11822
rect 3104 6462 3322 7170
rect 5250 6806 5444 6976
rect 14954 6414 15190 6542
rect 27126 6432 27316 6816
rect -390 4704 -180 4940
rect 30504 4716 30624 4900
rect 18236 3130 18560 3278
rect 24388 2334 24740 2774
rect -1394 1446 -862 1776
rect 3078 1672 3768 1912
rect 14938 1532 15204 1766
rect 26916 1602 27242 1842
rect 2094 598 2358 946
rect 18238 32 18554 206
rect 30738 -20 31282 142
<< metal2 >>
rect 12448 22430 12692 22480
rect 12448 22238 12484 22430
rect 12650 22238 12692 22430
rect 12448 22200 12692 22238
rect 15404 22428 15678 22480
rect 15404 22266 15448 22428
rect 15656 22266 15678 22428
rect 15404 22224 15678 22266
rect 30838 20854 31168 20898
rect -702 20774 186 20802
rect -1260 20566 -866 20608
rect -1260 20206 -1196 20566
rect -920 20206 -866 20566
rect -702 20596 -366 20774
rect 128 20596 186 20774
rect -702 20550 186 20596
rect -1260 20172 -866 20206
rect -700 5550 -564 20550
rect 30838 20530 30894 20854
rect 31122 20530 31168 20854
rect 30838 20466 31168 20530
rect 29714 20022 29936 20048
rect 29714 19740 29734 20022
rect 29898 19982 29936 20022
rect 29898 19897 30586 19982
rect 29898 19740 29936 19897
rect 29714 19708 29936 19740
rect 29614 13706 30026 13782
rect 28420 13470 29294 13556
rect 20550 13434 20722 13452
rect 7344 13398 7588 13414
rect 7344 13304 7372 13398
rect 7562 13304 7588 13398
rect 7344 13288 7588 13304
rect -432 12388 -148 12470
rect -432 12220 -416 12388
rect -200 12220 -148 12388
rect -700 5506 -490 5550
rect -700 5388 -670 5506
rect -698 5310 -670 5388
rect -524 5310 -490 5506
rect -698 5290 -490 5310
rect -432 4972 -148 12220
rect 7480 12292 7588 13288
rect 20550 13304 20574 13434
rect 20696 13304 20722 13434
rect 20550 13284 20722 13304
rect 20550 12292 20650 13284
rect 28420 13002 28550 13470
rect 29202 13002 29294 13470
rect 7480 12276 7760 12292
rect 7480 12192 7500 12276
rect 7740 12192 7760 12276
rect 7480 12180 7760 12192
rect 7488 12178 7760 12180
rect 20520 12274 20664 12292
rect 20520 12170 20544 12274
rect 20650 12170 20664 12274
rect 20520 12158 20664 12170
rect 28420 11822 29294 13002
rect 29614 12276 29684 13706
rect 29966 12276 30026 13706
rect 30501 13033 30586 19897
rect 29614 12216 30026 12276
rect 30500 12268 30586 13033
rect 28420 11662 28520 11822
rect 29240 11662 29294 11822
rect 28420 11606 29294 11662
rect 30271 12182 30586 12268
rect 30271 11335 30357 12182
rect 30888 12100 31102 20466
rect 30527 11998 31102 12100
rect 30527 11451 30629 11998
rect 30888 11996 31102 11998
rect 30696 11822 31318 11858
rect 30696 11570 30746 11822
rect 31286 11570 31318 11822
rect 30696 11538 31318 11570
rect 30527 11392 30901 11451
rect 30640 11349 30901 11392
rect 30271 11292 30500 11335
rect 30799 11312 30901 11349
rect 30271 11249 30586 11292
rect 30402 11118 30586 11249
rect 30799 11215 30904 11312
rect 3078 7170 3362 7220
rect 3078 6462 3104 7170
rect 3322 6618 3362 7170
rect 5210 6980 5476 7006
rect 5210 6850 5236 6980
rect 5376 6976 5476 6980
rect 5210 6806 5250 6850
rect 5444 6806 5476 6976
rect 5210 6782 5476 6806
rect 27076 6816 27366 6882
rect 3322 6462 3464 6618
rect 3078 6426 3464 6462
rect 14924 6542 15220 6562
rect 3078 6346 3462 6426
rect 14924 6414 14954 6542
rect 15190 6414 15220 6542
rect 27076 6510 27126 6816
rect 14924 6388 15220 6414
rect 26906 6432 27126 6510
rect 27316 6432 27366 6816
rect 26906 6396 27366 6432
rect -432 4940 -146 4972
rect -432 4704 -390 4940
rect -180 4704 -146 4940
rect -432 4670 -146 4704
rect 3284 1974 3462 6346
rect 3000 1912 3836 1974
rect -1442 1776 -820 1820
rect -1442 1446 -1394 1776
rect -862 1446 -820 1776
rect 3000 1672 3078 1912
rect 3768 1672 3836 1912
rect 14956 1798 15186 6388
rect 18200 3278 18582 3290
rect 18200 3130 18236 3278
rect 18560 3130 18582 3278
rect 3000 1618 3836 1672
rect 14916 1766 15230 1798
rect 14916 1532 14938 1766
rect 15204 1532 15230 1766
rect 14916 1500 15230 1532
rect -1442 1406 -820 1446
rect 2046 946 2394 988
rect 2046 598 2094 946
rect 2358 598 2394 946
rect 2046 558 2394 598
rect 18200 238 18582 3130
rect 24328 2774 24778 2802
rect 24328 2334 24388 2774
rect 24740 2334 24778 2774
rect 24328 2282 24778 2334
rect 26906 1878 27122 6396
rect 30500 4938 30586 11118
rect 30828 5836 30904 11215
rect 30716 5774 30974 5836
rect 30716 5280 30742 5774
rect 30930 5280 30974 5774
rect 30716 5240 30974 5280
rect 30474 4900 30656 4938
rect 30474 4716 30504 4900
rect 30624 4716 30656 4900
rect 30474 4676 30656 4716
rect 30500 4542 30586 4676
rect 26874 1842 27270 1878
rect 26874 1602 26916 1842
rect 27242 1602 27270 1842
rect 26874 1564 27270 1602
rect 18198 206 18582 238
rect 18198 32 18238 206
rect 18554 32 18582 206
rect 18198 0 18582 32
rect 30696 142 31318 170
rect 30696 -20 30738 142
rect 31282 -20 31318 142
rect 30696 -42 31318 -20
<< via2 >>
rect 12484 22238 12650 22430
rect 15448 22266 15656 22428
rect -1196 20206 -920 20566
rect -416 12220 -200 12388
rect -670 5310 -524 5506
rect 7500 12192 7740 12276
rect 20544 12170 20650 12274
rect 29684 12276 29966 13706
rect 30746 11570 31286 11822
rect 5236 6976 5376 6980
rect 5236 6850 5250 6976
rect 5250 6850 5376 6976
rect -1394 1446 -862 1776
rect 2094 598 2358 946
rect 24388 2334 24740 2774
rect 30742 5280 30930 5774
rect 30738 -20 31282 142
<< metal3 >>
rect 12448 22430 12692 22480
rect 12448 22238 12484 22430
rect 12650 22238 12692 22430
rect 12448 22200 12692 22238
rect 15404 22428 15678 22480
rect 15404 22266 15448 22428
rect 15656 22266 15678 22428
rect 15404 22224 15678 22266
rect -1260 20566 -866 20608
rect -1260 20206 -1196 20566
rect -920 20206 -866 20566
rect -1260 20172 -866 20206
rect 29614 13706 30026 13782
rect 29614 12436 29684 13706
rect -436 12388 3452 12428
rect -436 12220 -416 12388
rect -200 12220 3452 12388
rect 7488 12276 7760 12292
rect 7488 12254 7500 12276
rect -436 12194 3452 12220
rect 7480 12192 7500 12254
rect 7740 12252 7760 12276
rect 20520 12274 20664 12292
rect 20520 12252 20544 12274
rect 7740 12192 20544 12252
rect 7480 12182 20544 12192
rect 7480 12180 7760 12182
rect 7488 12178 7760 12180
rect 20520 12170 20544 12182
rect 20650 12170 20664 12274
rect 25176 12276 29684 12436
rect 29966 12276 30026 13706
rect 25176 12216 30026 12276
rect 20520 12158 20664 12170
rect 30696 11822 31318 11858
rect 30696 11570 30746 11822
rect 31286 11570 31318 11822
rect 30696 11538 31318 11570
rect 4738 7054 5412 7096
rect 4738 6844 4796 7054
rect 5348 6980 5412 7054
rect 5376 6914 5412 6980
rect 9666 7074 10122 7112
rect 5376 6850 6742 6914
rect 5348 6844 6742 6850
rect 4738 6828 6742 6844
rect 9666 6882 9742 7074
rect 10064 6882 10122 7074
rect 9666 6828 10122 6882
rect 20148 7088 20526 7130
rect 20148 6854 20176 7088
rect 20466 6854 20526 7088
rect 20148 6830 20526 6854
rect 25028 7078 25490 7124
rect 25028 6870 25100 7078
rect 25442 6870 25490 7078
rect 25028 6828 25490 6870
rect 4738 6810 5412 6828
rect 30716 5774 30974 5836
rect 14524 5552 14840 5590
rect -698 5548 -490 5550
rect -698 5506 1218 5548
rect -698 5310 -670 5506
rect -524 5310 1218 5506
rect -698 5290 1218 5310
rect 14524 5336 14570 5552
rect 14794 5336 14840 5552
rect 30716 5550 30742 5774
rect 14524 5298 14840 5336
rect 29896 5292 30742 5550
rect 30716 5280 30742 5292
rect 30930 5280 30974 5774
rect 30716 5240 30974 5280
rect 3708 3616 11106 3846
rect 19010 3614 25206 3848
rect 24328 2774 24778 2802
rect 24328 2334 24388 2774
rect 24740 2334 24778 2774
rect 24328 2282 24778 2334
rect -1442 1776 -820 1820
rect -1442 1446 -1394 1776
rect -862 1446 -820 1776
rect -1442 1406 -820 1446
rect 2046 946 2394 988
rect 2046 598 2094 946
rect 2358 598 2394 946
rect 2046 558 2394 598
rect 30696 142 31318 170
rect 30696 -20 30738 142
rect 31282 -20 31318 142
rect 30696 -42 31318 -20
<< via3 >>
rect 12484 22238 12650 22430
rect 15448 22266 15656 22428
rect -1196 20206 -920 20566
rect 30746 11570 31286 11822
rect 4796 6980 5348 7054
rect 4796 6850 5236 6980
rect 5236 6850 5348 6980
rect 4796 6844 5348 6850
rect 9742 6882 10064 7074
rect 20176 6854 20466 7088
rect 25100 6870 25442 7078
rect 14570 5336 14794 5552
rect 15728 5322 15974 5524
rect 24388 2334 24740 2774
rect -1394 1446 -862 1776
rect 2094 598 2358 946
rect 30738 -20 31282 142
<< metal4 >>
rect -1442 20566 -820 23352
rect 12448 22430 12692 22480
rect 12448 22238 12484 22430
rect 12650 22290 12692 22430
rect 15404 22428 15678 22480
rect 15404 22298 15448 22428
rect 12650 22238 13734 22290
rect 12448 22200 13734 22238
rect 14236 22266 15448 22298
rect 15656 22266 15678 22428
rect 14236 22224 15678 22266
rect 14236 22222 15510 22224
rect 12480 22194 13734 22200
rect 13646 21756 13732 22194
rect 13646 21750 13738 21756
rect 13646 21690 13836 21750
rect 13750 21460 13836 21690
rect -1442 20206 -1196 20566
rect -920 20206 -820 20566
rect 13647 21374 13836 21460
rect 13647 21372 13738 21374
rect 13647 20326 13731 21372
rect 14248 20396 14324 22222
rect 13647 20242 13982 20326
rect -1442 1776 -820 20206
rect 13866 20162 13982 20242
rect 13890 19954 13982 20162
rect 13866 17618 13982 19954
rect 13888 17406 13982 17618
rect 13866 17126 13982 17406
rect 13888 16914 13982 17126
rect 13866 15604 13982 16914
rect 13888 15392 13982 15604
rect 13866 12698 13982 15392
rect 13868 12576 13982 12698
rect 14132 20320 14324 20396
rect 13868 11464 13948 12576
rect 9600 11340 9782 11344
rect 13770 11340 13948 11464
rect 9600 11194 13948 11340
rect 14132 11296 14208 20320
rect 30696 11822 31318 23396
rect 30696 11570 30746 11822
rect 31286 11570 31318 11822
rect 14132 11220 20334 11296
rect 9600 7112 9782 11194
rect 20258 7130 20334 11220
rect 4686 7096 4922 7106
rect 4686 7054 5412 7096
rect 4686 6844 4796 7054
rect 5348 6844 5412 7054
rect 4686 6810 5412 6844
rect 9600 7074 10122 7112
rect 9600 6882 9742 7074
rect 10064 6882 10122 7074
rect 9600 6832 10122 6882
rect 9666 6828 10122 6832
rect 20148 7088 20526 7130
rect 20148 6854 20176 7088
rect 20466 6854 20526 7088
rect 25028 7078 25490 7124
rect 25028 7032 25100 7078
rect 20148 6830 20526 6854
rect 24452 6870 25100 7032
rect 25442 6870 25490 7078
rect 24452 6828 25490 6870
rect 4686 3292 4922 6810
rect 16184 6406 16564 6446
rect 2268 3274 4922 3292
rect -1442 1446 -1394 1776
rect -862 1446 -820 1776
rect -1442 -266 -820 1446
rect 2260 3106 4922 3274
rect 13852 5958 16584 6406
rect 2260 988 2412 3106
rect 2046 946 2412 988
rect 2046 598 2094 946
rect 2358 598 2412 946
rect 2046 588 2412 598
rect 2046 558 2394 588
rect 13852 -514 14260 5958
rect 14524 5552 14840 5590
rect 14524 5336 14570 5552
rect 14794 5336 14840 5552
rect 14524 5298 14840 5336
rect 14524 -520 14838 5298
rect 15168 -528 15482 5958
rect 15698 5524 16012 5544
rect 15698 5322 15728 5524
rect 15974 5322 16012 5524
rect 15698 -538 16012 5322
rect 16184 -542 16564 5958
rect 24452 2802 24644 6828
rect 24328 2774 24778 2802
rect 24328 2334 24388 2774
rect 24740 2334 24778 2774
rect 24328 2282 24778 2334
rect 30696 326 31318 11570
rect 30694 142 31318 326
rect 30694 -20 30738 142
rect 31282 -20 31318 142
rect 30694 -44 31318 -20
use analog_buffer  analog_buffer_0
timestamp 1717178954
transform -1 0 6842 0 1 4126
box -742 -726 6842 7776
use analog_buffer  analog_buffer_1
timestamp 1717178954
transform 1 0 23598 0 1 4126
box -742 -726 6842 7776
use analog_buffer  analog_buffer_2
timestamp 1717178954
transform 1 0 8216 0 1 4126
box -742 -726 6842 7776
use analog_buffer  analog_buffer_3
timestamp 1717178954
transform -1 0 21962 0 1 4126
box -742 -726 6842 7776
use current_source  current_source_0
timestamp 1717178954
transform -1 0 30384 0 -1 20752
box -54 544 936 8966
use filter22M  filter22M_0
timestamp 1717178954
transform -1 0 28160 0 1 12002
box -2 0 13828 11358
use filter22M  filter22M_1
timestamp 1717178954
transform 1 0 2 0 1 12000
box -2 0 13828 11358
use oscillator_20MHZ  oscillator_20MHZ_0
timestamp 1717178954
transform -1 0 29159 0 1 2
box 0 -2 26159 1646
use oscillator_21MHZ  oscillator_21MHZ_0
timestamp 1717178954
transform 1 0 6000 0 -1 3282
box 0 -1 18074 1646
<< labels >>
flabel metal4 -1442 1776 -820 23352 0 FreeSans 1600 0 0 0 VCC
port 7 nsew
flabel metal4 2268 3106 4922 3292 0 FreeSans 1600 0 0 0 OSCA
flabel metal4 24388 2334 24740 2774 0 FreeSans 1600 0 0 0 OSCB
flabel metal4 30696 142 31318 23396 0 FreeSans 1600 0 0 0 VSS
flabel metal3 29896 5292 30742 5550 0 FreeSans 1600 0 0 0 OSCB_BUF
flabel metal3 -524 5290 1218 5548 0 FreeSans 1600 0 0 0 OSCA_BUF
flabel metal4 9600 11194 13948 11340 0 FreeSans 1600 0 0 0 FIL_OUTA
flabel metal4 14132 11220 20334 11296 0 FreeSans 1600 0 0 0 FIL_OUTB
flabel metal4 14524 -520 14838 5336 0 FreeSans 1600 0 0 0 OUTA
port 8 nsew
flabel metal4 15698 -538 16012 5322 0 FreeSans 1600 0 0 0 OUTB
port 9 nsew
flabel metal4 30696 11822 31318 23396 0 FreeSans 1600 0 0 0 VSS
port 10 nsew
<< end >>
