magic
tech sky130A
magscale 1 2
timestamp 1716504190
<< pwell >>
rect -415 -2596 415 2596
<< psubdiff >>
rect -379 2526 -283 2560
rect 283 2526 379 2560
rect -379 2464 -345 2526
rect 345 2464 379 2526
rect -379 -2526 -345 -2464
rect 345 -2526 379 -2464
rect -379 -2560 -283 -2526
rect 283 -2560 379 -2526
<< psubdiffcont >>
rect -283 2526 283 2560
rect -379 -2464 -345 2464
rect 345 -2464 379 2464
rect -283 -2560 283 -2526
<< poly >>
rect -249 2414 -183 2430
rect -249 2380 -233 2414
rect -199 2380 -183 2414
rect -249 2000 -183 2380
rect -249 -2380 -183 -2000
rect -249 -2414 -233 -2380
rect -199 -2414 -183 -2380
rect -249 -2430 -183 -2414
rect -141 2414 -75 2430
rect -141 2380 -125 2414
rect -91 2380 -75 2414
rect -141 2000 -75 2380
rect -141 -2380 -75 -2000
rect -141 -2414 -125 -2380
rect -91 -2414 -75 -2380
rect -141 -2430 -75 -2414
rect -33 2414 33 2430
rect -33 2380 -17 2414
rect 17 2380 33 2414
rect -33 2000 33 2380
rect -33 -2380 33 -2000
rect -33 -2414 -17 -2380
rect 17 -2414 33 -2380
rect -33 -2430 33 -2414
rect 75 2414 141 2430
rect 75 2380 91 2414
rect 125 2380 141 2414
rect 75 2000 141 2380
rect 75 -2380 141 -2000
rect 75 -2414 91 -2380
rect 125 -2414 141 -2380
rect 75 -2430 141 -2414
rect 183 2414 249 2430
rect 183 2380 199 2414
rect 233 2380 249 2414
rect 183 2000 249 2380
rect 183 -2380 249 -2000
rect 183 -2414 199 -2380
rect 233 -2414 249 -2380
rect 183 -2430 249 -2414
<< polycont >>
rect -233 2380 -199 2414
rect -233 -2414 -199 -2380
rect -125 2380 -91 2414
rect -125 -2414 -91 -2380
rect -17 2380 17 2414
rect -17 -2414 17 -2380
rect 91 2380 125 2414
rect 91 -2414 125 -2380
rect 199 2380 233 2414
rect 199 -2414 233 -2380
<< npolyres >>
rect -249 -2000 -183 2000
rect -141 -2000 -75 2000
rect -33 -2000 33 2000
rect 75 -2000 141 2000
rect 183 -2000 249 2000
<< locali >>
rect -379 2526 -283 2560
rect 283 2526 379 2560
rect -379 2464 -345 2526
rect 345 2464 379 2526
rect -249 2380 -233 2414
rect -199 2380 -183 2414
rect -141 2380 -125 2414
rect -91 2380 -75 2414
rect -33 2380 -17 2414
rect 17 2380 33 2414
rect 75 2380 91 2414
rect 125 2380 141 2414
rect 183 2380 199 2414
rect 233 2380 249 2414
rect -249 -2414 -233 -2380
rect -199 -2414 -183 -2380
rect -141 -2414 -125 -2380
rect -91 -2414 -75 -2380
rect -33 -2414 -17 -2380
rect 17 -2414 33 -2380
rect 75 -2414 91 -2380
rect 125 -2414 141 -2380
rect 183 -2414 199 -2380
rect 233 -2414 249 -2380
rect -379 -2526 -345 -2464
rect 345 -2526 379 -2464
rect -379 -2560 -283 -2526
rect 283 -2560 379 -2526
<< viali >>
rect -233 2380 -199 2414
rect -125 2380 -91 2414
rect -17 2380 17 2414
rect 91 2380 125 2414
rect 199 2380 233 2414
rect -233 2017 -199 2380
rect -125 2017 -91 2380
rect -17 2017 17 2380
rect 91 2017 125 2380
rect 199 2017 233 2380
rect -233 -2380 -199 -2017
rect -125 -2380 -91 -2017
rect -17 -2380 17 -2017
rect 91 -2380 125 -2017
rect 199 -2380 233 -2017
rect -233 -2414 -199 -2380
rect -125 -2414 -91 -2380
rect -17 -2414 17 -2380
rect 91 -2414 125 -2380
rect 199 -2414 233 -2380
<< metal1 >>
rect -239 2414 -193 2426
rect -239 2017 -233 2414
rect -199 2017 -193 2414
rect -239 2005 -193 2017
rect -131 2414 -85 2426
rect -131 2017 -125 2414
rect -91 2017 -85 2414
rect -131 2005 -85 2017
rect -23 2414 23 2426
rect -23 2017 -17 2414
rect 17 2017 23 2414
rect -23 2005 23 2017
rect 85 2414 131 2426
rect 85 2017 91 2414
rect 125 2017 131 2414
rect 85 2005 131 2017
rect 193 2414 239 2426
rect 193 2017 199 2414
rect 233 2017 239 2414
rect 193 2005 239 2017
rect -239 -2017 -193 -2005
rect -239 -2414 -233 -2017
rect -199 -2414 -193 -2017
rect -239 -2426 -193 -2414
rect -131 -2017 -85 -2005
rect -131 -2414 -125 -2017
rect -91 -2414 -85 -2017
rect -131 -2426 -85 -2414
rect -23 -2017 23 -2005
rect -23 -2414 -17 -2017
rect 17 -2414 23 -2017
rect -23 -2426 23 -2414
rect 85 -2017 131 -2005
rect 85 -2414 91 -2017
rect 125 -2414 131 -2017
rect 85 -2426 131 -2414
rect 193 -2017 239 -2005
rect 193 -2414 199 -2017
rect 233 -2414 239 -2017
rect 193 -2426 239 -2414
<< properties >>
string FIXED_BBOX -362 -2543 362 2543
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.330 l 20 m 1 nx 5 wmin 0.330 lmin 1.650 rho 48.2 val 2.921k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
