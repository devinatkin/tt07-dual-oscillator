magic
tech sky130A
magscale 1 2
timestamp 1716498465
<< nwell >>
rect 5222 480 8676 1260
rect 8650 478 8676 480
<< pwell >>
rect 3866 2450 8675 5872
rect 3868 1262 8675 2450
rect 4360 1261 8675 1262
<< metal1 >>
rect 3498 5694 4066 5808
rect 7983 5710 8423 5713
rect 3868 4114 4066 5694
rect 6968 5690 7175 5698
rect 7451 5690 7658 5710
rect 7983 5695 8473 5710
rect 6612 5687 7658 5690
rect 5026 5671 5129 5675
rect 4773 5660 4969 5667
rect 4367 5641 4969 5660
rect 4314 5566 4969 5641
rect 4314 4678 4432 5566
rect 4842 4678 4969 5566
rect 4314 4568 4969 4678
rect 5026 5552 5348 5671
rect 5026 5250 5129 5552
rect 5279 5250 5348 5552
rect 5026 5177 5348 5250
rect 5512 5667 5719 5679
rect 5926 5667 6133 5683
rect 5512 5572 6133 5667
rect 5512 5236 5614 5572
rect 5994 5236 6133 5572
rect 5026 5143 5340 5177
rect 4314 4545 4961 4568
rect 5026 4545 5129 5143
rect 5512 5136 6133 5236
rect 5512 5135 5876 5136
rect 4451 4541 4961 4545
rect 5512 4541 5719 5135
rect 5988 4545 6133 5136
rect 6493 5518 7658 5687
rect 6493 4549 6700 5518
rect 6968 4560 7175 5518
rect 7451 4572 7658 5518
rect 7945 5572 8473 5695
rect 7945 5142 8082 5572
rect 8360 5142 8473 5572
rect 7945 5043 8473 5142
rect 7945 4557 8152 5043
rect 3797 4002 4066 4114
rect 1838 3925 4066 4002
rect 3797 3868 4066 3925
rect 3262 3127 3427 3156
rect 3262 2843 3289 3127
rect 3405 2843 3427 3127
rect 3262 2796 3427 2843
rect 2021 2613 2034 2708
rect 2189 2613 2199 2708
rect 2021 2589 2199 2613
rect 1580 2346 1851 2377
rect 1580 2190 1619 2346
rect 1800 2190 1851 2346
rect 1580 2154 1851 2190
rect 3868 1222 4066 3868
rect 5208 1080 5480 1261
rect 3200 947 3467 976
rect 3200 776 3233 947
rect 3427 776 3467 947
rect 3200 754 3467 776
rect 5314 360 5480 1080
rect 1298 -2523 1471 -646
rect 5425 -834 5725 -799
rect 5425 -1018 5446 -834
rect 5692 -1018 5725 -834
rect 5425 -1035 5725 -1018
rect 4789 -1197 5681 -1173
rect 4789 -1318 4825 -1197
rect 4989 -1318 5681 -1197
rect 4789 -1347 5681 -1318
rect 3449 -2122 3642 -2113
rect 1638 -2199 3643 -2122
rect 1638 -2200 3468 -2199
rect 3449 -2325 3468 -2200
rect 3630 -2200 3643 -2199
rect 3630 -2325 3642 -2200
rect 3449 -2345 3642 -2325
rect 3774 -2518 3976 -2506
rect 3534 -2592 3976 -2518
rect 3534 -2604 3930 -2592
rect 5143 -2604 5444 -2532
<< via1 >>
rect 3289 2843 3405 3127
rect 2034 2613 2189 2711
rect 1619 2190 1800 2346
rect 3233 776 3427 947
rect 5446 -1018 5692 -834
rect 4825 -1318 4989 -1197
rect 3468 -2325 3630 -2199
rect 4126 -2481 4178 -2223
<< metal2 >>
rect 3286 3158 3433 3773
rect 3170 3127 3433 3158
rect 3170 2843 3289 3127
rect 3405 3117 3433 3127
rect 3405 2843 3432 3117
rect 2021 2711 2199 2720
rect 2021 2613 2034 2711
rect 2189 2613 2199 2711
rect 1580 2346 1851 2377
rect 1580 2190 1619 2346
rect 1800 2190 1851 2346
rect 1580 2154 1851 2190
rect 2021 1978 2199 2613
rect 3170 2294 3432 2843
rect 3780 2609 4167 2610
rect 3780 2568 4249 2609
rect 3170 2166 3710 2294
rect 3170 2164 3432 2166
rect 2021 1673 2043 1978
rect 2170 1673 2199 1978
rect 2021 1642 2199 1673
rect 3596 1440 3710 2166
rect 3780 1758 3827 2568
rect 4160 1758 4249 2568
rect 3780 1716 4249 1758
rect 3780 1700 4365 1716
rect 3596 1212 3614 1440
rect 3684 1212 3710 1440
rect 4106 1381 4365 1700
rect 5534 1506 5850 1575
rect 5534 1462 6091 1506
rect 4682 1416 5194 1454
rect 3200 951 3467 976
rect 3200 947 3300 951
rect 3200 776 3233 947
rect 3441 820 3467 951
rect 3427 776 3467 820
rect 3200 754 3467 776
rect 3596 528 3710 1212
rect 3596 486 3779 528
rect 3596 273 3629 486
rect 3731 273 3779 486
rect 3596 236 3779 273
rect 2763 -294 2937 -283
rect 2763 -385 2784 -294
rect 2924 -385 2937 -294
rect 2763 -1097 2937 -385
rect 3599 -873 3779 236
rect 4107 -512 4249 1381
rect 4682 1258 4736 1416
rect 5112 1258 5194 1416
rect 4682 756 5194 1258
rect 5534 1244 5603 1462
rect 5535 1178 5603 1244
rect 6033 1178 6091 1462
rect 5535 1135 6091 1178
rect 5535 587 5800 1135
rect 4662 534 4936 556
rect 4662 329 4698 534
rect 4906 329 4936 534
rect 4662 -429 4936 329
rect 5535 340 5577 587
rect 5767 340 5800 587
rect 5535 316 5800 340
rect 4107 -710 4134 -512
rect 4224 -710 4249 -512
rect 4107 -752 4249 -710
rect 3599 -995 3618 -873
rect 3759 -995 3779 -873
rect 3599 -1009 3779 -995
rect 5425 -834 5725 -799
rect 5425 -1018 5446 -834
rect 5692 -1018 5725 -834
rect 5425 -1035 5725 -1018
rect 2763 -1259 2778 -1097
rect 2911 -1259 2937 -1097
rect 2763 -1268 2937 -1259
rect 4786 -1197 5035 -1173
rect 4786 -1318 4825 -1197
rect 4989 -1318 5035 -1197
rect 3447 -2199 3741 -2121
rect 3447 -2325 3468 -2199
rect 3630 -2202 3741 -2199
rect 3447 -2402 3469 -2325
rect 3709 -2402 3741 -2202
rect 3447 -2415 3741 -2402
rect 4062 -2203 4270 -2190
rect 4062 -2397 4076 -2203
rect 4252 -2397 4270 -2203
rect 4062 -2481 4126 -2397
rect 4178 -2481 4270 -2397
rect 4786 -2201 5035 -1318
rect 4786 -2392 4816 -2201
rect 5001 -2392 5035 -2201
rect 4786 -2418 5035 -2392
rect 4062 -2506 4270 -2481
<< via2 >>
rect 1619 2190 1800 2346
rect 2043 1673 2170 1978
rect 3827 1758 4160 2568
rect 3614 1212 3684 1440
rect 3300 947 3441 951
rect 3300 820 3427 947
rect 3427 820 3441 947
rect 3629 273 3731 486
rect 2784 -385 2924 -294
rect 4736 1258 5112 1416
rect 5603 1178 6033 1462
rect 4698 329 4906 534
rect 5577 340 5767 587
rect 4134 -710 4224 -512
rect 3618 -995 3759 -873
rect 5446 -1018 5692 -834
rect 2778 -1259 2911 -1097
rect 3469 -2325 3630 -2202
rect 3630 -2325 3709 -2202
rect 3469 -2402 3709 -2325
rect 4076 -2223 4252 -2203
rect 4076 -2397 4126 -2223
rect 4126 -2397 4178 -2223
rect 4178 -2397 4252 -2223
rect 4816 -2392 5001 -2201
<< metal3 >>
rect 3780 2572 4286 2619
rect 1580 2346 1851 2377
rect 1580 2190 1619 2346
rect 1800 2190 1851 2346
rect 1580 2154 1851 2190
rect 3780 1751 3809 2572
rect 4165 1751 4286 2572
rect 3780 1700 4286 1751
rect 5536 1462 6091 1506
rect 3566 1440 5195 1455
rect 3566 1212 3614 1440
rect 3684 1416 5195 1440
rect 3684 1258 4736 1416
rect 5112 1258 5195 1416
rect 3684 1212 5195 1258
rect 3566 1200 5195 1212
rect 5536 1178 5603 1462
rect 6033 1178 6091 1462
rect 5536 1135 6091 1178
rect 3266 951 3533 1018
rect 3266 820 3300 951
rect 3441 820 3533 951
rect 3266 796 3533 820
rect 4665 587 5793 621
rect 4665 534 5577 587
rect 2423 486 3757 509
rect 2423 273 3629 486
rect 3731 273 3757 486
rect 4665 329 4698 534
rect 4906 340 5577 534
rect 5767 340 5793 587
rect 4906 329 5793 340
rect 4665 312 5793 329
rect 2423 235 3757 273
rect 4097 -512 5699 -479
rect 4097 -710 4134 -512
rect 4224 -710 5699 -512
rect 4097 -751 5699 -710
rect 7758 -734 7962 -482
rect 5414 -834 5714 -818
rect 5414 -851 5446 -834
rect 3599 -873 5446 -851
rect 3599 -995 3618 -873
rect 3759 -995 5446 -873
rect 3599 -1009 5446 -995
rect 5414 -1018 5446 -1009
rect 5692 -1018 5714 -834
rect 5414 -1054 5714 -1018
rect 3447 -2201 5032 -2185
rect 3447 -2202 4816 -2201
rect 3447 -2402 3469 -2202
rect 3709 -2203 4816 -2202
rect 3709 -2397 4076 -2203
rect 4252 -2392 4816 -2203
rect 5001 -2392 5032 -2201
rect 4252 -2397 5032 -2392
rect 3709 -2402 5032 -2397
rect 3447 -2416 5032 -2402
<< via3 >>
rect 3809 2568 4165 2572
rect 3809 1758 3827 2568
rect 3827 1758 4160 2568
rect 4160 1758 4165 2568
rect 3809 1751 4165 1758
rect 5603 1178 6033 1462
<< metal4 >>
rect 4173 2611 4304 4315
rect 3771 2572 4304 2611
rect 3771 1751 3809 2572
rect 4165 1751 4304 2572
rect 3771 1716 4304 1751
rect 3771 1700 4277 1716
rect 5536 1462 6094 1878
rect 5536 1178 5603 1462
rect 6033 1178 6094 1462
rect 5536 1135 6094 1178
use active-resistor  active-resistor_0
timestamp 1716495568
transform 1 0 418 0 1 -844
box 3450 -1784 4804 2106
use activeload  activeload_0
timestamp 1716496561
transform 1 0 1092 0 1 2452
box 0 0 2774 3420
use indiff  indiff_0
timestamp 1716478495
transform 1 0 1524 0 1 -480
box -382 -304 2344 2930
use second_stage  second_stage_0
timestamp 1716496561
transform 1 0 5450 0 1 -2466
box -228 -164 3226 2946
use sky130_fd_pr__cap_mim_m3_1_NY928X  sky130_fd_pr__cap_mim_m3_1_NY928X_0
timestamp 1716478495
transform -1 0 6394 0 -1 2980
box -2186 -1340 2186 1340
use tail_current  tail_current_0
timestamp 1716495288
transform 1 0 1092 0 1 -2628
box 0 0 2774 1844
<< labels >>
flabel metal1 1638 -2200 3643 -2122 0 FreeSans 800 0 0 0 IBIAS
port 0 nsew
flabel metal3 3441 796 3533 1018 0 FreeSans 800 0 0 0 INB
port 1 nsew
flabel metal3 1800 2154 1851 2377 0 FreeSans 800 0 0 0 INA
port 2 nsew
flabel space 3508 -2592 4000 -2506 0 FreeSans 640 0 0 0 VSS
port 3 nsew
flabel metal1 3820 5694 4038 5808 0 FreeSans 640 0 0 0 VCC
port 4 nsew
flabel metal3 7758 -734 7962 -482 0 FreeSans 640 0 0 0 OUT
port 5 nsew
flabel metal1 3534 -2604 3930 -2518 0 FreeSans 320 0 0 0 VSS
port 6 nsew
<< end >>
