magic
tech sky130A
magscale 1 2
timestamp 1716523272
<< nwell >>
rect 3450 2006 4804 2104
rect 3450 1934 3582 2006
rect 3450 1754 3478 1934
rect 3524 1918 3582 1934
rect 3816 1918 4804 2006
rect 3524 1754 4804 1918
rect 3450 418 4804 1754
rect 3450 411 3616 418
rect 3806 411 4804 418
rect 3450 360 3597 411
rect 3820 360 4804 411
rect 3450 359 3616 360
rect 3806 359 4804 360
rect 3450 281 3540 359
rect 3814 348 4804 359
rect 4084 288 4804 348
rect 3814 281 4804 288
rect 3450 264 3616 281
rect 3806 264 4804 281
rect 3450 188 4804 264
rect 3450 128 3612 188
rect 3634 173 4804 188
rect 3450 61 3634 128
rect 3796 61 4804 173
rect 3450 -364 4804 61
<< pwell >>
rect 3450 -478 4804 -364
rect 3450 -562 3822 -478
rect 3848 -520 4804 -478
rect 3848 -560 3874 -520
rect 3926 -560 4804 -520
rect 3450 -576 3848 -562
rect 3958 -576 4804 -560
rect 3450 -588 3874 -576
rect 3926 -588 4804 -576
rect 3450 -1574 4804 -588
rect 3450 -1684 3606 -1574
rect 3640 -1684 4804 -1574
rect 3450 -1784 4804 -1684
<< viali >>
rect 3582 2036 3810 2070
rect 4056 1936 4284 1970
rect 4442 1936 4670 1970
rect 3486 1778 3520 1892
rect 3872 1606 3906 1834
rect 3872 450 3906 1440
rect 3960 450 3994 1440
rect 3486 -806 3520 -678
rect 3486 -1042 3520 -914
rect 3486 -1322 3520 -1194
rect 3486 -1652 3520 -1524
rect 3582 -1748 3910 -1714
<< metal1 >>
rect 3450 2070 4804 2104
rect 3450 2036 3582 2070
rect 3810 2036 4804 2070
rect 3450 2006 4804 2036
rect 3450 1892 3582 2006
rect 3816 1970 4804 2006
rect 3450 1778 3486 1892
rect 3520 1778 3634 1892
rect 3450 1736 3634 1778
rect 3692 1886 3760 1968
rect 3816 1936 4056 1970
rect 4284 1936 4442 1970
rect 4670 1936 4804 1970
rect 3816 1924 4804 1936
rect 3692 1772 3796 1886
rect 3754 418 3796 1772
rect 3858 1834 3928 1924
rect 3858 1606 3872 1834
rect 3906 1606 3928 1834
rect 4120 1826 4606 1884
rect 4066 1776 4134 1780
rect 3858 1522 3928 1606
rect 4002 1766 4134 1776
rect 4002 1604 4014 1766
rect 4098 1604 4134 1766
rect 4002 1594 4134 1604
rect 3858 1440 4008 1522
rect 3858 450 3872 1440
rect 3906 450 3960 1440
rect 3994 450 4008 1440
rect 3858 398 4008 450
rect 3752 346 3798 397
rect 4066 386 4134 1594
rect 4226 730 4498 1790
rect 4600 1776 4668 1780
rect 4596 1768 4708 1776
rect 4596 1606 4610 1768
rect 4694 1606 4708 1768
rect 4596 1594 4708 1606
rect 4226 426 4268 730
rect 4450 426 4498 730
rect 4226 382 4498 426
rect 4600 386 4668 1594
rect 3713 345 3798 346
rect 3570 342 3798 345
rect 3570 330 3731 342
rect 3739 330 3798 342
rect 3570 299 3798 330
rect 3570 264 3616 299
rect 4084 290 4606 348
rect 4084 288 4328 290
rect 3570 188 3622 264
rect 4084 238 4144 288
rect 3752 204 4144 238
rect 3570 -140 3612 188
rect 3752 173 3954 204
rect 3650 95 3954 173
rect 3752 -184 3954 95
rect 3646 -242 3954 -184
rect 3904 -476 3952 -242
rect 3468 -678 3636 -570
rect 3468 -806 3486 -678
rect 3520 -806 3636 -678
rect 3468 -914 3636 -806
rect 3468 -1042 3486 -914
rect 3520 -1042 3636 -914
rect 3468 -1194 3636 -1042
rect 3468 -1322 3486 -1194
rect 3520 -1322 3636 -1194
rect 3468 -1524 3636 -1322
rect 3468 -1652 3486 -1524
rect 3520 -1574 3636 -1524
rect 3520 -1652 3606 -1574
rect 3702 -1650 3770 -500
rect 3904 -520 3964 -476
rect 3926 -573 3964 -520
rect 3856 -588 3874 -576
rect 3898 -588 3964 -573
rect 3856 -616 3964 -588
rect 3856 -1580 3952 -616
rect 3468 -1684 3606 -1652
rect 3468 -1688 3636 -1684
rect 3468 -1714 4776 -1688
rect 3468 -1748 3582 -1714
rect 3910 -1748 4776 -1714
rect 3468 -1760 4776 -1748
<< via1 >>
rect 4014 1604 4098 1766
rect 4610 1606 4694 1768
rect 4268 426 4450 730
<< metal2 >>
rect 4002 1768 4708 1776
rect 4002 1766 4610 1768
rect 4002 1604 4014 1766
rect 4098 1606 4610 1766
rect 4694 1606 4708 1768
rect 4098 1604 4708 1606
rect 4002 1594 4708 1604
rect 4228 730 4492 766
rect 4228 426 4268 730
rect 4450 426 4492 730
rect 4228 398 4492 426
use sky130_fd_pr__nfet_01v8_VNG24X  sky130_fd_pr__nfet_01v8_VNG24X_0
timestamp 1716523272
transform 1 0 3747 0 1 -1074
box -296 -710 296 710
use sky130_fd_pr__pfet_01v8_lvt_B5E2Q5  sky130_fd_pr__pfet_01v8_lvt_B5E2Q5_0
timestamp 1716523272
transform 1 0 3696 0 1 -45
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_lvt_E4WS6L  sky130_fd_pr__pfet_01v8_lvt_E4WS6L_0
timestamp 1716523272
transform 1 0 4557 0 1 1088
box -246 -919 246 919
use sky130_fd_pr__pfet_01v8_lvt_EG9S6L  sky130_fd_pr__pfet_01v8_lvt_EG9S6L_0
timestamp 1716523272
transform 1 0 4171 0 1 1088
box -246 -919 246 919
use sky130_fd_pr__pfet_01v8_lvt_NZC8UH  sky130_fd_pr__pfet_01v8_lvt_NZC8UH_0
timestamp 1716523272
transform 1 0 3696 0 1 1137
box -246 -969 246 969
<< labels >>
flabel metal1 3702 -1650 3770 -500 0 FreeSans 320 0 0 0 IBIAS
port 7 nsew
flabel metal1 3816 1924 4056 2104 0 FreeSans 320 0 0 0 VCC
port 8 nsew
flabel metal1 3910 -1760 4776 -1688 0 FreeSans 320 0 0 0 VSS
port 9 nsew
flabel metal2 4098 1594 4610 1776 0 FreeSans 320 0 0 0 RP
port 10 nsew
flabel via1 4268 426 4450 730 0 FreeSans 320 0 0 0 RN
port 11 nsew
flabel metal1 3904 -520 3952 -184 0 FreeSans 320 0 0 0 Rbias
<< end >>
