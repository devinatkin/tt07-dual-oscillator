magic
tech sky130A
magscale 1 2
timestamp 1716335449
<< nwell >>
rect -246 -1955 246 1955
<< pmoslvt >>
rect -50 736 50 1736
rect -50 -500 50 500
rect -50 -1736 50 -736
<< pdiff >>
rect -108 1724 -50 1736
rect -108 748 -96 1724
rect -62 748 -50 1724
rect -108 736 -50 748
rect 50 1724 108 1736
rect 50 748 62 1724
rect 96 748 108 1724
rect 50 736 108 748
rect -108 488 -50 500
rect -108 -488 -96 488
rect -62 -488 -50 488
rect -108 -500 -50 -488
rect 50 488 108 500
rect 50 -488 62 488
rect 96 -488 108 488
rect 50 -500 108 -488
rect -108 -748 -50 -736
rect -108 -1724 -96 -748
rect -62 -1724 -50 -748
rect -108 -1736 -50 -1724
rect 50 -748 108 -736
rect 50 -1724 62 -748
rect 96 -1724 108 -748
rect 50 -1736 108 -1724
<< pdiffc >>
rect -96 748 -62 1724
rect 62 748 96 1724
rect -96 -488 -62 488
rect 62 -488 96 488
rect -96 -1724 -62 -748
rect 62 -1724 96 -748
<< nsubdiff >>
rect -210 1885 -114 1919
rect 114 1885 210 1919
rect -210 1823 -176 1885
rect 176 1823 210 1885
rect -210 -1885 -176 -1823
rect 176 -1885 210 -1823
rect -210 -1919 -114 -1885
rect 114 -1919 210 -1885
<< nsubdiffcont >>
rect -114 1885 114 1919
rect -210 -1823 -176 1823
rect 176 -1823 210 1823
rect -114 -1919 114 -1885
<< poly >>
rect -50 1817 50 1833
rect -50 1783 -34 1817
rect 34 1783 50 1817
rect -50 1736 50 1783
rect -50 689 50 736
rect -50 655 -34 689
rect 34 655 50 689
rect -50 639 50 655
rect -50 581 50 597
rect -50 547 -34 581
rect 34 547 50 581
rect -50 500 50 547
rect -50 -547 50 -500
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect -50 -597 50 -581
rect -50 -655 50 -639
rect -50 -689 -34 -655
rect 34 -689 50 -655
rect -50 -736 50 -689
rect -50 -1783 50 -1736
rect -50 -1817 -34 -1783
rect 34 -1817 50 -1783
rect -50 -1833 50 -1817
<< polycont >>
rect -34 1783 34 1817
rect -34 655 34 689
rect -34 547 34 581
rect -34 -581 34 -547
rect -34 -689 34 -655
rect -34 -1817 34 -1783
<< locali >>
rect -210 1885 -114 1919
rect 114 1885 210 1919
rect -210 1823 -176 1885
rect 176 1823 210 1885
rect -50 1783 -34 1817
rect 34 1783 50 1817
rect -96 1724 -62 1740
rect -96 732 -62 748
rect 62 1724 96 1740
rect 62 732 96 748
rect -50 655 -34 689
rect 34 655 50 689
rect -50 547 -34 581
rect 34 547 50 581
rect -96 488 -62 504
rect -96 -504 -62 -488
rect 62 488 96 504
rect 62 -504 96 -488
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect -50 -689 -34 -655
rect 34 -689 50 -655
rect -96 -748 -62 -732
rect -96 -1740 -62 -1724
rect 62 -748 96 -732
rect 62 -1740 96 -1724
rect -50 -1817 -34 -1783
rect 34 -1817 50 -1783
rect -210 -1885 -176 -1823
rect 176 -1885 210 -1823
rect -210 -1919 -114 -1885
rect 114 -1919 210 -1885
<< viali >>
rect -34 1783 34 1817
rect -96 748 -62 1724
rect 62 748 96 1724
rect -34 655 34 689
rect -34 547 34 581
rect -96 -488 -62 488
rect 62 -488 96 488
rect -34 -581 34 -547
rect -34 -689 34 -655
rect -96 -1724 -62 -748
rect 62 -1724 96 -748
rect -34 -1817 34 -1783
<< metal1 >>
rect -46 1817 46 1823
rect -46 1783 -34 1817
rect 34 1783 46 1817
rect -46 1777 46 1783
rect -102 1724 -56 1736
rect -102 748 -96 1724
rect -62 748 -56 1724
rect -102 736 -56 748
rect 56 1724 102 1736
rect 56 748 62 1724
rect 96 748 102 1724
rect 56 736 102 748
rect -46 689 46 695
rect -46 655 -34 689
rect 34 655 46 689
rect -46 649 46 655
rect -46 581 46 587
rect -46 547 -34 581
rect 34 547 46 581
rect -46 541 46 547
rect -102 488 -56 500
rect -102 -488 -96 488
rect -62 -488 -56 488
rect -102 -500 -56 -488
rect 56 488 102 500
rect 56 -488 62 488
rect 96 -488 102 488
rect 56 -500 102 -488
rect -46 -547 46 -541
rect -46 -581 -34 -547
rect 34 -581 46 -547
rect -46 -587 46 -581
rect -46 -655 46 -649
rect -46 -689 -34 -655
rect 34 -689 46 -655
rect -46 -695 46 -689
rect -102 -748 -56 -736
rect -102 -1724 -96 -748
rect -62 -1724 -56 -748
rect -102 -1736 -56 -1724
rect 56 -748 102 -736
rect 56 -1724 62 -748
rect 96 -1724 102 -748
rect 56 -1736 102 -1724
rect -46 -1783 46 -1777
rect -46 -1817 -34 -1783
rect 34 -1817 46 -1783
rect -46 -1823 46 -1817
<< properties >>
string FIXED_BBOX -193 -1902 193 1902
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5.0 l 0.5 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
