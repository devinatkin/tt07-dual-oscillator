magic
tech sky130A
magscale 1 2
timestamp 1717035347
<< pwell >>
rect -216 -3596 216 3596
<< psubdiff >>
rect -180 3526 -84 3560
rect 84 3526 180 3560
rect -180 3464 -146 3526
rect 146 3464 180 3526
rect -180 -3526 -146 -3464
rect 146 -3526 180 -3464
rect -180 -3560 -84 -3526
rect 84 -3560 180 -3526
<< psubdiffcont >>
rect -84 3526 84 3560
rect -180 -3464 -146 3464
rect 146 -3464 180 3464
rect -84 -3560 84 -3526
<< poly >>
rect -50 3414 50 3430
rect -50 3380 -34 3414
rect 34 3380 50 3414
rect -50 3000 50 3380
rect -50 -3380 50 -3000
rect -50 -3414 -34 -3380
rect 34 -3414 50 -3380
rect -50 -3430 50 -3414
<< polycont >>
rect -34 3380 34 3414
rect -34 -3414 34 -3380
<< npolyres >>
rect -50 -3000 50 3000
<< locali >>
rect -180 3526 -84 3560
rect 84 3526 180 3560
rect -180 3464 -146 3526
rect 146 3464 180 3526
rect -50 3380 -34 3414
rect 34 3380 50 3414
rect -50 -3414 -34 -3380
rect 34 -3414 50 -3380
rect -180 -3526 -146 -3464
rect 146 -3526 180 -3464
rect -180 -3560 -84 -3526
rect 84 -3560 180 -3526
<< viali >>
rect -34 3380 34 3414
rect -34 3017 34 3380
rect -34 -3380 34 -3017
rect -34 -3414 34 -3380
<< metal1 >>
rect -40 3414 40 3426
rect -40 3017 -34 3414
rect 34 3017 40 3414
rect -40 3005 40 3017
rect -40 -3017 40 -3005
rect -40 -3414 -34 -3017
rect 34 -3414 40 -3017
rect -40 -3426 40 -3414
<< properties >>
string FIXED_BBOX -163 -3543 163 3543
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.5 l 30 m 1 nx 1 wmin 0.330 lmin 1.650 rho 48.2 val 2.892k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
