magic
tech sky130A
timestamp 1716523272
<< pwell >>
rect 0 0 1387 922
<< psubdiff >>
rect 46 849 156 866
rect 1150 849 1360 866
rect 46 810 63 849
rect 46 43 63 79
rect 1343 813 1360 849
rect 1343 43 1360 82
rect 46 26 237 43
rect 1231 26 1360 43
<< psubdiffcont >>
rect 156 849 1150 866
rect 46 79 63 810
rect 1343 82 1360 813
rect 237 26 1231 43
<< locali >>
rect 46 849 156 866
rect 1150 849 1360 866
rect 46 810 63 849
rect 46 43 63 79
rect 1343 813 1360 849
rect 1343 43 1360 82
rect 46 26 237 43
rect 1231 26 1360 43
<< viali >>
rect 237 26 1208 43
<< metal1 >>
rect 273 812 1274 816
rect 273 788 693 812
rect 688 786 693 788
rect 729 788 1274 812
rect 729 786 733 788
rect 688 779 733 786
rect 240 766 282 772
rect 498 766 540 772
rect 757 768 795 772
rect 240 689 246 766
rect 272 689 282 766
rect 240 680 282 689
rect 247 270 270 680
rect 376 380 399 766
rect 498 684 503 766
rect 533 684 540 766
rect 498 680 540 684
rect 356 368 423 380
rect 356 279 363 368
rect 411 279 423 368
rect 356 270 423 279
rect 505 271 528 680
rect 633 372 656 767
rect 757 684 762 768
rect 792 684 795 768
rect 1013 767 1050 772
rect 757 679 795 684
rect 626 366 665 372
rect 626 286 632 366
rect 659 286 665 366
rect 626 278 665 286
rect 633 271 656 278
rect 763 271 786 679
rect 891 372 914 767
rect 1013 687 1018 767
rect 1044 687 1050 767
rect 1013 680 1050 687
rect 882 367 920 372
rect 882 283 888 367
rect 915 283 920 367
rect 882 277 920 283
rect 891 271 914 277
rect 1020 271 1043 680
rect 1150 372 1173 767
rect 1274 766 1306 773
rect 1274 685 1278 766
rect 1304 685 1306 766
rect 1274 680 1306 685
rect 1142 367 1182 372
rect 1142 282 1148 367
rect 1176 282 1182 367
rect 1142 277 1182 282
rect 1150 271 1173 277
rect 688 259 733 261
rect 688 253 692 259
rect 273 233 692 253
rect 728 253 733 259
rect 728 233 1274 253
rect 273 228 1274 233
rect 356 69 422 78
rect 356 61 365 69
rect 46 43 365 61
rect 413 61 422 69
rect 413 43 1360 61
rect 46 26 237 43
rect 1208 26 1360 43
rect 46 18 1360 26
<< via1 >>
rect 693 786 729 812
rect 246 689 272 766
rect 503 684 533 766
rect 363 279 411 368
rect 762 684 792 768
rect 632 286 659 366
rect 1018 687 1044 767
rect 888 283 915 367
rect 1278 685 1304 766
rect 1148 282 1176 367
rect 692 233 728 259
rect 365 43 413 69
rect 365 30 413 43
<< metal2 >>
rect 688 812 733 816
rect 688 786 693 812
rect 729 786 733 812
rect 240 768 282 772
rect 240 685 246 768
rect 277 685 282 768
rect 240 680 282 685
rect 498 766 540 772
rect 498 683 503 766
rect 534 683 540 766
rect 498 680 540 683
rect 356 368 423 380
rect 356 279 363 368
rect 411 279 423 368
rect 356 270 423 279
rect 622 368 668 375
rect 622 282 628 368
rect 662 282 668 368
rect 622 274 668 282
rect 356 69 422 270
rect 688 259 733 786
rect 756 768 799 773
rect 756 683 762 768
rect 792 766 799 768
rect 793 683 799 766
rect 756 679 799 683
rect 1013 767 1050 772
rect 1013 688 1017 767
rect 1046 688 1050 767
rect 1013 687 1018 688
rect 1044 687 1050 688
rect 1013 680 1050 687
rect 1270 766 1307 773
rect 1270 765 1278 766
rect 1304 765 1307 766
rect 1270 684 1275 765
rect 1306 684 1307 765
rect 1270 679 1307 684
rect 878 368 924 374
rect 878 283 886 368
rect 916 283 924 368
rect 878 274 924 283
rect 1140 367 1183 372
rect 1140 282 1142 367
rect 1178 282 1183 367
rect 1140 277 1183 282
rect 688 233 692 259
rect 728 233 733 259
rect 688 228 733 233
rect 356 30 365 69
rect 413 30 422 69
rect 356 18 422 30
<< via2 >>
rect 246 766 277 768
rect 246 689 272 766
rect 272 689 277 766
rect 246 685 277 689
rect 503 684 533 766
rect 533 684 534 766
rect 503 683 534 684
rect 369 280 406 365
rect 628 366 662 368
rect 628 286 632 366
rect 632 286 659 366
rect 659 286 662 366
rect 628 282 662 286
rect 762 684 792 766
rect 792 684 793 766
rect 762 683 793 684
rect 1017 688 1018 767
rect 1018 688 1044 767
rect 1044 688 1046 767
rect 1275 685 1278 765
rect 1278 685 1304 765
rect 1304 685 1306 765
rect 1275 684 1306 685
rect 886 367 916 368
rect 886 283 888 367
rect 888 283 915 367
rect 915 283 916 367
rect 1142 282 1148 367
rect 1148 282 1176 367
rect 1176 282 1178 367
<< metal3 >>
rect 1111 772 1333 773
rect 243 768 1333 772
rect 243 685 246 768
rect 277 767 1333 768
rect 277 766 1017 767
rect 277 685 503 766
rect 243 683 503 685
rect 534 683 762 766
rect 793 688 1017 766
rect 1046 765 1333 767
rect 1046 688 1275 765
rect 793 684 1275 688
rect 1306 684 1333 765
rect 793 683 1333 684
rect 243 680 1333 683
rect 363 370 416 375
rect 623 370 669 376
rect 877 370 927 377
rect 1134 370 1356 371
rect 247 368 1356 370
rect 247 365 628 368
rect 247 280 369 365
rect 406 282 628 365
rect 662 283 886 368
rect 916 367 1356 368
rect 916 283 1142 367
rect 662 282 1142 283
rect 1178 282 1356 367
rect 406 280 1356 282
rect 247 278 1356 280
rect 363 269 416 278
rect 623 274 669 278
rect 877 273 927 278
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_1
timestamp 1716523272
transform 1 0 323 0 1 522
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_2
timestamp 1716523272
transform 1 0 452 0 1 522
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_3
timestamp 1716523272
transform 1 0 1097 0 1 522
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_4
timestamp 1716523272
transform 1 0 581 0 1 522
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_5
timestamp 1716523272
transform 1 0 710 0 1 522
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_6
timestamp 1716523272
transform 1 0 839 0 1 522
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_7
timestamp 1716523272
transform 1 0 968 0 1 522
box -79 -294 79 294
use sky130_fd_pr__nfet_01v8_U654K6  sky130_fd_pr__nfet_01v8_U654K6_8
timestamp 1716523272
transform 1 0 1226 0 1 522
box -79 -294 79 294
<< labels >>
flabel pwell 46 18 1360 61 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 728 228 1274 253 0 FreeSans 400 0 0 0 IBIAS
port 4 nsew
flabel metal3 277 680 503 772 0 FreeSans 400 0 0 0 TAILV
port 5 nsew
flabel pwell 78 18 591 57 0 FreeSans 320 0 0 0 VSS
port 6 nsew
<< end >>
