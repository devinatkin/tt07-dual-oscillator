magic
tech sky130A
timestamp 1717178954
<< metal3 >>
rect -247 4640 2817 4670
rect -247 3127 -215 4640
rect -165 4563 2736 4593
rect -165 3893 -127 4563
rect 2706 3896 2736 4563
rect 2782 3928 2817 4640
rect -165 3847 -160 3893
rect -128 3847 -126 3893
rect 2706 3891 2749 3896
rect -165 3844 -126 3847
rect 1231 3853 1268 3857
rect -165 3837 -127 3844
rect -165 3130 -130 3837
rect 1231 3813 1234 3853
rect 1266 3813 1268 3853
rect -247 3123 -195 3127
rect -247 3085 -243 3123
rect -200 3085 -195 3123
rect -247 2362 -195 3085
rect -247 2324 -244 2362
rect -201 2324 -195 2362
rect -247 2116 -195 2324
rect -247 2078 -242 2116
rect -199 2078 -195 2116
rect -247 2073 -195 2078
rect -165 3067 -129 3130
rect -165 2368 -127 3067
rect -165 2121 -123 2368
rect -247 1499 -216 2073
rect -247 846 -217 1499
rect -165 1466 -121 2121
rect -171 1389 -121 1466
rect -171 878 -129 1389
rect -164 877 -129 878
rect -164 847 -121 877
rect -164 846 -120 847
rect -247 842 -195 846
rect -247 804 -245 842
rect -202 804 -195 842
rect -247 784 -195 804
rect -165 800 -119 846
rect -247 -180 -208 784
rect -165 749 -120 800
rect -176 745 -120 749
rect -176 699 -131 745
rect -176 82 -135 699
rect 1231 662 1268 3813
rect 2706 3850 2714 3891
rect 2746 3850 2749 3891
rect 2706 3842 2749 3850
rect 1309 3089 1346 3095
rect 1309 3050 1311 3089
rect 1343 3050 1346 3089
rect 2706 3072 2736 3842
rect 2786 3838 2817 3928
rect 2782 3127 2817 3838
rect 2769 3124 2817 3127
rect 2769 3085 2772 3124
rect 2812 3085 2817 3124
rect 2769 3081 2817 3085
rect 2706 3053 2740 3072
rect 1309 2326 1346 3050
rect 2704 3042 2740 3053
rect 2704 2996 2734 3042
rect 2704 2966 2736 2996
rect 2706 2680 2736 2966
rect 2706 2650 2737 2680
rect 1309 2289 1311 2326
rect 1345 2289 1346 2326
rect 1309 2153 1346 2289
rect 1309 2116 1311 2153
rect 1345 2116 1346 2153
rect 1309 1457 1346 2116
rect 2707 2312 2737 2650
rect 2776 2364 2817 3081
rect 2811 2325 2817 2364
rect 2776 2321 2817 2325
rect 2707 2282 2739 2312
rect -176 41 -175 82
rect -136 41 -135 82
rect -176 38 -135 41
rect 1229 629 1268 662
rect 1229 589 1234 629
rect 1266 589 1268 629
rect 1229 155 1268 589
rect 1229 44 1233 155
rect 1265 44 1268 155
rect 1229 40 1268 44
rect 1308 1395 1347 1457
rect 1308 1394 1348 1395
rect 1308 1357 1311 1394
rect 1345 1357 1348 1394
rect 1308 1354 1348 1357
rect 1308 155 1347 1354
rect 2707 759 2737 2282
rect 2785 2121 2817 2321
rect 2767 2118 2817 2121
rect 2767 2079 2771 2118
rect 2811 2079 2817 2118
rect 2767 2075 2817 2079
rect 2785 847 2817 2075
rect 2767 843 2817 847
rect 2767 804 2771 843
rect 2811 804 2817 843
rect 2767 800 2817 804
rect 2707 722 2755 759
rect 1308 44 1312 155
rect 1344 44 1347 155
rect 2725 94 2755 722
rect 1308 40 1347 44
rect 2701 89 2755 94
rect 2701 43 2707 89
rect 2752 43 2755 89
rect 2701 39 2755 43
rect -176 37 -129 38
rect -172 -75 -129 37
rect -172 -104 -128 -75
rect 2725 -93 2755 39
rect 1398 -104 1448 -100
rect -172 -120 -127 -104
rect 1398 -120 1403 -104
rect -172 -146 1403 -120
rect 1444 -116 1448 -104
rect 1444 -120 1599 -116
rect 2724 -120 2755 -93
rect 1444 -146 2755 -120
rect -172 -150 1459 -146
rect 1573 -150 2755 -146
rect 1503 -177 1547 -176
rect 1503 -180 1506 -177
rect -247 -209 1506 -180
rect 1544 -180 1547 -177
rect 2787 -180 2817 800
rect 1544 -209 2817 -180
rect -247 -210 2817 -209
<< via3 >>
rect -160 3847 -128 3893
rect 1234 3813 1266 3853
rect -243 3085 -200 3123
rect -244 2324 -201 2362
rect -242 2078 -199 2116
rect -245 804 -202 842
rect 2714 3850 2746 3891
rect 1311 3050 1343 3089
rect 2772 3085 2812 3124
rect 1311 2289 1345 2326
rect 1311 2116 1345 2153
rect 2776 2325 2811 2364
rect -175 41 -136 82
rect 1234 589 1266 629
rect 1233 44 1265 155
rect 1311 1357 1345 1394
rect 2771 2079 2811 2118
rect 2771 804 2811 843
rect 1312 44 1344 155
rect 2707 43 2752 89
rect 1403 -146 1444 -104
rect 1506 -209 1544 -177
<< metal4 >>
rect -165 3896 -99 3897
rect 41 3896 1004 4403
rect -165 3893 1004 3896
rect -165 3847 -160 3893
rect -128 3847 1004 3893
rect 1585 3896 2547 4404
rect 1585 3891 2749 3896
rect -165 3842 1004 3847
rect 41 3840 1004 3842
rect 1139 3853 1453 3857
rect 1139 3813 1234 3853
rect 1266 3813 1453 3853
rect 1585 3850 2714 3891
rect 2746 3850 2749 3891
rect 1585 3842 2749 3850
rect 1139 3809 1453 3813
rect 41 3127 1003 3643
rect -247 3123 1003 3127
rect -247 3085 -243 3123
rect -200 3085 1003 3123
rect 1585 3127 2547 3643
rect 1585 3124 2817 3127
rect 1309 3089 1346 3090
rect -247 3081 1003 3085
rect 1137 3050 1311 3089
rect 1343 3050 1450 3089
rect 1585 3085 2772 3124
rect 2812 3085 2817 3124
rect 1585 3081 2817 3085
rect 1137 3049 1450 3050
rect 40 2366 1002 2882
rect -247 2362 1002 2366
rect -247 2324 -244 2362
rect -201 2324 1002 2362
rect 1585 2367 2547 2883
rect 1585 2351 2586 2367
rect 2707 2364 2817 2367
rect 2707 2351 2776 2364
rect -247 2320 1002 2324
rect 1137 2326 1450 2327
rect 1137 2289 1311 2326
rect 1345 2289 1450 2326
rect 1585 2325 2776 2351
rect 2811 2325 2817 2364
rect 1585 2321 2817 2325
rect 1137 2287 1450 2289
rect 1136 2153 1451 2154
rect 39 2120 1001 2121
rect -247 2116 1001 2120
rect -247 2078 -242 2116
rect -199 2078 1001 2116
rect 1136 2116 1311 2153
rect 1345 2116 1451 2153
rect 1136 2114 1451 2116
rect 1586 2121 2548 2122
rect 1586 2118 2818 2121
rect -247 2074 1001 2078
rect 39 1559 1001 2074
rect 1586 2079 2771 2118
rect 2811 2079 2818 2118
rect 1586 2075 2818 2079
rect 1586 1560 2548 2075
rect 1136 1394 1451 1395
rect 39 846 1001 1361
rect 1136 1357 1311 1394
rect 1345 1357 1451 1394
rect 1136 1355 1451 1357
rect -248 842 1001 846
rect -248 804 -245 842
rect -202 804 1001 842
rect -248 800 1001 804
rect 1585 847 2547 1362
rect 1585 843 2817 847
rect 1585 804 2771 843
rect 2811 804 2817 843
rect 1585 801 2817 804
rect 1585 800 2547 801
rect 39 799 1001 800
rect 1136 629 1450 634
rect 39 93 1001 601
rect 1136 589 1234 629
rect 1266 589 1450 629
rect 1136 586 1450 589
rect -178 82 1001 93
rect -178 41 -175 82
rect -136 41 1001 82
rect -178 39 1001 41
rect 1229 155 1268 158
rect 1229 44 1233 155
rect 1265 44 1268 155
rect -178 38 -71 39
rect 1229 -205 1268 44
rect 1308 155 1347 158
rect 1308 44 1312 155
rect 1344 44 1347 155
rect 1308 -205 1347 44
rect 1585 93 2547 601
rect 1585 69 2586 93
rect 2701 89 2755 93
rect 2701 69 2707 89
rect 1585 43 2707 69
rect 2752 43 2755 89
rect 1585 39 2755 43
rect 1398 -104 1448 -94
rect 1398 -146 1403 -104
rect 1444 -146 1448 -104
rect 1398 -206 1448 -146
rect 1503 -177 1553 -154
rect 1503 -209 1506 -177
rect 1544 -209 1553 -177
rect 1503 -210 1553 -209
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_0
timestamp 1717178954
transform 1 0 593 0 1 1080
box -593 -320 593 320
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_1
timestamp 1717178954
transform -1 0 1993 0 -1 1081
box -593 -320 593 320
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_2
timestamp 1717178954
transform 1 0 596 0 1 4123
box -593 -320 593 320
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_3
timestamp 1717178954
transform 1 0 593 0 1 1840
box -593 -320 593 320
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_4
timestamp 1717178954
transform 1 0 594 0 1 2601
box -593 -320 593 320
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_5
timestamp 1717178954
transform 1 0 595 0 1 3362
box -593 -320 593 320
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_6
timestamp 1717178954
transform 1 0 593 0 1 320
box -593 -320 593 320
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_7
timestamp 1717178954
transform -1 0 1993 0 -1 320
box -593 -320 593 320
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_8
timestamp 1717178954
transform -1 0 1993 0 -1 4123
box -593 -320 593 320
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_9
timestamp 1717178954
transform -1 0 1994 0 -1 1841
box -593 -320 593 320
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_10
timestamp 1717178954
transform -1 0 1993 0 -1 2602
box -593 -320 593 320
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_11
timestamp 1717178954
transform -1 0 1993 0 -1 3362
box -593 -320 593 320
<< labels >>
flabel metal4 1229 -205 1268 44 0 FreeSans 80 0 0 0 CAPA_N
port 1 nsew
flabel metal4 1308 -205 1347 44 0 FreeSans 80 0 0 0 CAPB_N
port 2 nsew
flabel metal4 1398 -206 1448 -100 0 FreeSans 80 0 0 0 CAPA_P
port 3 nsew
flabel metal4 1503 -160 1553 -154 0 FreeSans 80 0 0 0 CAPB_P
port 4 nsew
<< end >>
